magic
tech sky130A
magscale 1 2
timestamp 1641099986
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 251174 700992 251180 701004
rect 202840 700964 251180 700992
rect 202840 700952 202846 700964
rect 251174 700952 251180 700964
rect 251232 700952 251238 701004
rect 248322 700884 248328 700936
rect 248380 700924 248386 700936
rect 348786 700924 348792 700936
rect 248380 700896 348792 700924
rect 248380 700884 248386 700896
rect 348786 700884 348792 700896
rect 348844 700884 348850 700936
rect 154114 700816 154120 700868
rect 154172 700856 154178 700868
rect 255314 700856 255320 700868
rect 154172 700828 255320 700856
rect 154172 700816 154178 700828
rect 255314 700816 255320 700828
rect 255372 700816 255378 700868
rect 137830 700748 137836 700800
rect 137888 700788 137894 700800
rect 253934 700788 253940 700800
rect 137888 700760 253940 700788
rect 137888 700748 137894 700760
rect 253934 700748 253940 700760
rect 253992 700748 253998 700800
rect 245562 700680 245568 700732
rect 245620 700720 245626 700732
rect 413646 700720 413652 700732
rect 245620 700692 413652 700720
rect 245620 700680 245626 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 256786 700652 256792 700664
rect 89220 700624 256792 700652
rect 89220 700612 89226 700624
rect 256786 700612 256792 700624
rect 256844 700612 256850 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 256694 700584 256700 700596
rect 73028 700556 256700 700584
rect 73028 700544 73034 700556
rect 256694 700544 256700 700556
rect 256752 700544 256758 700596
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 41322 700516 41328 700528
rect 40552 700488 41328 700516
rect 40552 700476 40558 700488
rect 41322 700476 41328 700488
rect 41380 700476 41386 700528
rect 242802 700476 242808 700528
rect 242860 700516 242866 700528
rect 478506 700516 478512 700528
rect 242860 700488 478512 700516
rect 242860 700476 242866 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 24302 700408 24308 700460
rect 24360 700448 24366 700460
rect 259546 700448 259552 700460
rect 24360 700420 259552 700448
rect 24360 700408 24366 700420
rect 259546 700408 259552 700420
rect 259604 700408 259610 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 259454 700380 259460 700392
rect 8168 700352 259460 700380
rect 8168 700340 8174 700352
rect 259454 700340 259460 700352
rect 259512 700340 259518 700392
rect 295978 700340 295984 700392
rect 296036 700380 296042 700392
rect 300118 700380 300124 700392
rect 296036 700352 300124 700380
rect 296036 700340 296042 700352
rect 300118 700340 300124 700352
rect 300176 700340 300182 700392
rect 241330 700272 241336 700324
rect 241388 700312 241394 700324
rect 543458 700312 543464 700324
rect 241388 700284 543464 700312
rect 241388 700272 241394 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 218974 700204 218980 700256
rect 219032 700244 219038 700256
rect 252554 700244 252560 700256
rect 219032 700216 252560 700244
rect 219032 700204 219038 700216
rect 252554 700204 252560 700216
rect 252612 700204 252618 700256
rect 251082 700136 251088 700188
rect 251140 700176 251146 700188
rect 283834 700176 283840 700188
rect 251140 700148 283840 700176
rect 251140 700136 251146 700148
rect 283834 700136 283840 700148
rect 283892 700136 283898 700188
rect 249702 700068 249708 700120
rect 249760 700108 249766 700120
rect 267642 700108 267648 700120
rect 249760 700080 267648 700108
rect 249760 700068 249766 700080
rect 267642 700068 267648 700080
rect 267700 700068 267706 700120
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 233142 699660 233148 699712
rect 233200 699700 233206 699712
rect 235166 699700 235172 699712
rect 233200 699672 235172 699700
rect 233200 699660 233206 699672
rect 235166 699660 235172 699672
rect 235224 699660 235230 699712
rect 359458 699660 359464 699712
rect 359516 699700 359522 699712
rect 364978 699700 364984 699712
rect 359516 699672 364984 699700
rect 359516 699660 359522 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 461578 699660 461584 699712
rect 461636 699700 461642 699712
rect 462314 699700 462320 699712
rect 461636 699672 462320 699700
rect 461636 699660 461642 699672
rect 462314 699660 462320 699672
rect 462372 699660 462378 699712
rect 526438 699660 526444 699712
rect 526496 699700 526502 699712
rect 527174 699700 527180 699712
rect 526496 699672 527180 699700
rect 526496 699660 526502 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 237282 696940 237288 696992
rect 237340 696980 237346 696992
rect 580166 696980 580172 696992
rect 237340 696952 580172 696980
rect 237340 696940 237346 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 260834 683244 260840 683256
rect 3476 683216 260840 683244
rect 3476 683204 3482 683216
rect 260834 683204 260840 683216
rect 260892 683204 260898 683256
rect 238570 683136 238576 683188
rect 238628 683176 238634 683188
rect 580166 683176 580172 683188
rect 238628 683148 580172 683176
rect 238628 683136 238634 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 670760 3424 670812
rect 3476 670800 3482 670812
rect 262214 670800 262220 670812
rect 3476 670772 262220 670800
rect 3476 670760 3482 670772
rect 262214 670760 262220 670772
rect 262272 670760 262278 670812
rect 235902 670692 235908 670744
rect 235960 670732 235966 670744
rect 580166 670732 580172 670744
rect 235960 670704 580172 670732
rect 235960 670692 235966 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 262306 656928 262312 656940
rect 3476 656900 262312 656928
rect 3476 656888 3482 656900
rect 262306 656888 262312 656900
rect 262364 656888 262370 656940
rect 234522 643084 234528 643136
rect 234580 643124 234586 643136
rect 580166 643124 580172 643136
rect 234580 643096 580172 643124
rect 234580 643084 234586 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 263594 632108 263600 632120
rect 3476 632080 263600 632108
rect 3476 632068 3482 632080
rect 263594 632068 263600 632080
rect 263652 632068 263658 632120
rect 235810 630640 235816 630692
rect 235868 630680 235874 630692
rect 580166 630680 580172 630692
rect 235868 630652 580172 630680
rect 235868 630640 235874 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 264974 618304 264980 618316
rect 3200 618276 264980 618304
rect 3200 618264 3206 618276
rect 264974 618264 264980 618276
rect 265032 618264 265038 618316
rect 234430 616836 234436 616888
rect 234488 616876 234494 616888
rect 580166 616876 580172 616888
rect 234488 616848 580172 616876
rect 234488 616836 234494 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 263686 605860 263692 605872
rect 3292 605832 263692 605860
rect 3292 605820 3298 605832
rect 263686 605820 263692 605832
rect 263744 605820 263750 605872
rect 231670 590656 231676 590708
rect 231728 590696 231734 590708
rect 579798 590696 579804 590708
rect 231728 590668 579804 590696
rect 231728 590656 231734 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 371694 585352 371700 585404
rect 371752 585392 371758 585404
rect 513558 585392 513564 585404
rect 371752 585364 513564 585392
rect 371752 585352 371758 585364
rect 513558 585352 513564 585364
rect 513616 585352 513622 585404
rect 446398 585284 446404 585336
rect 446456 585324 446462 585336
rect 513374 585324 513380 585336
rect 446456 585296 513380 585324
rect 446456 585284 446462 585296
rect 513374 585284 513380 585296
rect 513432 585284 513438 585336
rect 425698 585216 425704 585268
rect 425756 585256 425762 585268
rect 516410 585256 516416 585268
rect 425756 585228 516416 585256
rect 425756 585216 425762 585228
rect 516410 585216 516416 585228
rect 516468 585216 516474 585268
rect 489178 584468 489184 584520
rect 489236 584508 489242 584520
rect 513926 584508 513932 584520
rect 489236 584480 513932 584508
rect 489236 584468 489242 584480
rect 513926 584468 513932 584480
rect 513984 584468 513990 584520
rect 485038 584400 485044 584452
rect 485096 584440 485102 584452
rect 513558 584440 513564 584452
rect 485096 584412 513564 584440
rect 485096 584400 485102 584412
rect 513558 584400 513564 584412
rect 513616 584400 513622 584452
rect 371786 584332 371792 584384
rect 371844 584372 371850 584384
rect 513742 584372 513748 584384
rect 371844 584344 513748 584372
rect 371844 584332 371850 584344
rect 513742 584332 513748 584344
rect 513800 584332 513806 584384
rect 500218 584264 500224 584316
rect 500276 584304 500282 584316
rect 516318 584304 516324 584316
rect 500276 584276 516324 584304
rect 500276 584264 500282 584276
rect 516318 584264 516324 584276
rect 516376 584264 516382 584316
rect 493318 584196 493324 584248
rect 493376 584236 493382 584248
rect 513834 584236 513840 584248
rect 493376 584208 513840 584236
rect 493376 584196 493382 584208
rect 513834 584196 513840 584208
rect 513892 584196 513898 584248
rect 490558 584128 490564 584180
rect 490616 584168 490622 584180
rect 513650 584168 513656 584180
rect 490616 584140 513656 584168
rect 490616 584128 490622 584140
rect 513650 584128 513656 584140
rect 513708 584128 513714 584180
rect 483658 584060 483664 584112
rect 483716 584100 483722 584112
rect 513374 584100 513380 584112
rect 483716 584072 513380 584100
rect 483716 584060 483722 584072
rect 513374 584060 513380 584072
rect 513432 584060 513438 584112
rect 430574 583992 430580 584044
rect 430632 584032 430638 584044
rect 516226 584032 516232 584044
rect 430632 584004 516232 584032
rect 430632 583992 430638 584004
rect 516226 583992 516232 584004
rect 516284 583992 516290 584044
rect 427814 583924 427820 583976
rect 427872 583964 427878 583976
rect 513282 583964 513288 583976
rect 427872 583936 513288 583964
rect 427872 583924 427878 583936
rect 513282 583924 513288 583936
rect 513340 583924 513346 583976
rect 444742 583856 444748 583908
rect 444800 583896 444806 583908
rect 447778 583896 447784 583908
rect 444800 583868 447784 583896
rect 444800 583856 444806 583868
rect 447778 583856 447784 583868
rect 447836 583856 447842 583908
rect 497458 583856 497464 583908
rect 497516 583896 497522 583908
rect 513466 583896 513472 583908
rect 497516 583868 513472 583896
rect 497516 583856 497522 583868
rect 513466 583856 513472 583868
rect 513524 583856 513530 583908
rect 516134 583720 516140 583772
rect 516192 583760 516198 583772
rect 524414 583760 524420 583772
rect 516192 583732 524420 583760
rect 516192 583720 516198 583732
rect 524414 583720 524420 583732
rect 524472 583720 524478 583772
rect 371602 581068 371608 581120
rect 371660 581108 371666 581120
rect 373994 581108 374000 581120
rect 371660 581080 374000 581108
rect 371660 581068 371666 581080
rect 373994 581068 374000 581080
rect 374052 581068 374058 581120
rect 371326 581000 371332 581052
rect 371384 581040 371390 581052
rect 378226 581040 378232 581052
rect 371384 581012 378232 581040
rect 371384 581000 371390 581012
rect 378226 581000 378232 581012
rect 378284 581000 378290 581052
rect 378778 580252 378784 580304
rect 378836 580292 378842 580304
rect 427814 580292 427820 580304
rect 378836 580264 427820 580292
rect 378836 580252 378842 580264
rect 427814 580252 427820 580264
rect 427872 580252 427878 580304
rect 371510 579776 371516 579828
rect 371568 579816 371574 579828
rect 377030 579816 377036 579828
rect 371568 579788 377036 579816
rect 371568 579776 371574 579788
rect 377030 579776 377036 579788
rect 377088 579776 377094 579828
rect 371602 579708 371608 579760
rect 371660 579748 371666 579760
rect 378778 579748 378784 579760
rect 371660 579720 378784 579748
rect 371660 579708 371666 579720
rect 378778 579708 378784 579720
rect 378836 579708 378842 579760
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 266354 579680 266360 579692
rect 3384 579652 266360 579680
rect 3384 579640 3390 579652
rect 266354 579640 266360 579652
rect 266412 579640 266418 579692
rect 371694 579640 371700 579692
rect 371752 579680 371758 579692
rect 380158 579680 380164 579692
rect 371752 579652 380164 579680
rect 371752 579640 371758 579652
rect 380158 579640 380164 579652
rect 380216 579640 380222 579692
rect 444742 579640 444748 579692
rect 444800 579680 444806 579692
rect 447870 579680 447876 579692
rect 444800 579652 447876 579680
rect 444800 579640 444806 579652
rect 447870 579640 447876 579652
rect 447928 579640 447934 579692
rect 444926 578416 444932 578468
rect 444984 578456 444990 578468
rect 448146 578456 448152 578468
rect 444984 578428 448152 578456
rect 444984 578416 444990 578428
rect 448146 578416 448152 578428
rect 448204 578416 448210 578468
rect 371326 578280 371332 578332
rect 371384 578320 371390 578332
rect 375466 578320 375472 578332
rect 371384 578292 375472 578320
rect 371384 578280 371390 578292
rect 375466 578280 375472 578292
rect 375524 578280 375530 578332
rect 371694 578212 371700 578264
rect 371752 578252 371758 578264
rect 379146 578252 379152 578264
rect 371752 578224 379152 578252
rect 371752 578212 371758 578224
rect 379146 578212 379152 578224
rect 379204 578212 379210 578264
rect 371234 578076 371240 578128
rect 371292 578116 371298 578128
rect 371786 578116 371792 578128
rect 371292 578088 371792 578116
rect 371292 578076 371298 578088
rect 371786 578076 371792 578088
rect 371844 578076 371850 578128
rect 378134 577464 378140 577516
rect 378192 577504 378198 577516
rect 430574 577504 430580 577516
rect 378192 577476 430580 577504
rect 378192 577464 378198 577476
rect 430574 577464 430580 577476
rect 430632 577464 430638 577516
rect 371418 576988 371424 577040
rect 371476 577028 371482 577040
rect 376754 577028 376760 577040
rect 371476 577000 376760 577028
rect 371476 576988 371482 577000
rect 376754 576988 376760 577000
rect 376812 576988 376818 577040
rect 371602 576920 371608 576972
rect 371660 576960 371666 576972
rect 378134 576960 378140 576972
rect 371660 576932 378140 576960
rect 371660 576920 371666 576932
rect 378134 576920 378140 576932
rect 378192 576920 378198 576972
rect 371694 576852 371700 576904
rect 371752 576892 371758 576904
rect 379054 576892 379060 576904
rect 371752 576864 379060 576892
rect 371752 576852 371758 576864
rect 379054 576852 379060 576864
rect 379112 576852 379118 576904
rect 371602 576104 371608 576156
rect 371660 576144 371666 576156
rect 425698 576144 425704 576156
rect 371660 576116 425704 576144
rect 371660 576104 371666 576116
rect 425698 576104 425704 576116
rect 425756 576104 425762 576156
rect 371694 575492 371700 575544
rect 371752 575532 371758 575544
rect 376938 575532 376944 575544
rect 371752 575504 376944 575532
rect 371752 575492 371758 575504
rect 376938 575492 376944 575504
rect 376996 575492 377002 575544
rect 444742 575492 444748 575544
rect 444800 575532 444806 575544
rect 448238 575532 448244 575544
rect 444800 575504 448244 575532
rect 444800 575492 444806 575504
rect 448238 575492 448244 575504
rect 448296 575492 448302 575544
rect 444558 574064 444564 574116
rect 444616 574104 444622 574116
rect 447962 574104 447968 574116
rect 444616 574076 447968 574104
rect 444616 574064 444622 574076
rect 447962 574064 447968 574076
rect 448020 574064 448026 574116
rect 371602 571480 371608 571532
rect 371660 571520 371666 571532
rect 375374 571520 375380 571532
rect 371660 571492 375380 571520
rect 371660 571480 371666 571492
rect 375374 571480 375380 571492
rect 375432 571480 375438 571532
rect 444834 571480 444840 571532
rect 444892 571520 444898 571532
rect 448054 571520 448060 571532
rect 444892 571492 448060 571520
rect 444892 571480 444898 571492
rect 448054 571480 448060 571492
rect 448112 571480 448118 571532
rect 371510 570256 371516 570308
rect 371568 570296 371574 570308
rect 376202 570296 376208 570308
rect 371568 570268 376208 570296
rect 371568 570256 371574 570268
rect 376202 570256 376208 570268
rect 376260 570256 376266 570308
rect 371602 569984 371608 570036
rect 371660 570024 371666 570036
rect 376018 570024 376024 570036
rect 371660 569996 376024 570024
rect 371660 569984 371666 569996
rect 376018 569984 376024 569996
rect 376076 569984 376082 570036
rect 371694 569916 371700 569968
rect 371752 569956 371758 569968
rect 376846 569956 376852 569968
rect 371752 569928 376852 569956
rect 371752 569916 371758 569928
rect 376846 569916 376852 569928
rect 376904 569916 376910 569968
rect 516134 568896 516140 568948
rect 516192 568936 516198 568948
rect 520366 568936 520372 568948
rect 516192 568908 520372 568936
rect 516192 568896 516198 568908
rect 520366 568896 520372 568908
rect 520424 568896 520430 568948
rect 444926 568556 444932 568608
rect 444984 568596 444990 568608
rect 449158 568596 449164 568608
rect 444984 568568 449164 568596
rect 444984 568556 444990 568568
rect 449158 568556 449164 568568
rect 449216 568556 449222 568608
rect 516226 568556 516232 568608
rect 516284 568596 516290 568608
rect 524598 568596 524604 568608
rect 516284 568568 524604 568596
rect 516284 568556 516290 568568
rect 524598 568556 524604 568568
rect 524656 568556 524662 568608
rect 516502 568012 516508 568064
rect 516560 568052 516566 568064
rect 516778 568052 516784 568064
rect 516560 568024 516784 568052
rect 516560 568012 516566 568024
rect 516778 568012 516784 568024
rect 516836 568012 516842 568064
rect 371510 567876 371516 567928
rect 371568 567916 371574 567928
rect 372982 567916 372988 567928
rect 371568 567888 372988 567916
rect 371568 567876 371574 567888
rect 372982 567876 372988 567888
rect 373040 567876 373046 567928
rect 371510 567740 371516 567792
rect 371568 567780 371574 567792
rect 371694 567780 371700 567792
rect 371568 567752 371700 567780
rect 371568 567740 371574 567752
rect 371694 567740 371700 567752
rect 371752 567740 371758 567792
rect 371602 567672 371608 567724
rect 371660 567712 371666 567724
rect 374638 567712 374644 567724
rect 371660 567684 374644 567712
rect 371660 567672 371666 567684
rect 374638 567672 374644 567684
rect 374696 567672 374702 567724
rect 516226 567332 516232 567384
rect 516284 567372 516290 567384
rect 521746 567372 521752 567384
rect 516284 567344 521752 567372
rect 516284 567332 516290 567344
rect 521746 567332 521752 567344
rect 521804 567332 521810 567384
rect 516134 567264 516140 567316
rect 516192 567304 516198 567316
rect 519354 567304 519360 567316
rect 516192 567276 519360 567304
rect 516192 567264 516198 567276
rect 519354 567264 519360 567276
rect 519412 567264 519418 567316
rect 516226 567196 516232 567248
rect 516284 567236 516290 567248
rect 516870 567236 516876 567248
rect 516284 567208 516876 567236
rect 516284 567196 516290 567208
rect 516870 567196 516876 567208
rect 516928 567196 516934 567248
rect 516594 567128 516600 567180
rect 516652 567128 516658 567180
rect 516612 567100 516640 567128
rect 516870 567100 516876 567112
rect 516612 567072 516876 567100
rect 516870 567060 516876 567072
rect 516928 567060 516934 567112
rect 516502 566992 516508 567044
rect 516560 567032 516566 567044
rect 516778 567032 516784 567044
rect 516560 567004 516784 567032
rect 516560 566992 516566 567004
rect 516778 566992 516784 567004
rect 516836 566992 516842 567044
rect 371786 566176 371792 566228
rect 371844 566216 371850 566228
rect 374178 566216 374184 566228
rect 371844 566188 374184 566216
rect 371844 566176 371850 566188
rect 374178 566176 374184 566188
rect 374236 566176 374242 566228
rect 516502 566040 516508 566092
rect 516560 566080 516566 566092
rect 520458 566080 520464 566092
rect 516560 566052 520464 566080
rect 516560 566040 516566 566052
rect 520458 566040 520464 566052
rect 520516 566040 520522 566092
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 267734 565876 267740 565888
rect 3476 565848 267740 565876
rect 3476 565836 3482 565848
rect 267734 565836 267740 565848
rect 267792 565836 267798 565888
rect 371786 565836 371792 565888
rect 371844 565876 371850 565888
rect 373258 565876 373264 565888
rect 371844 565848 373264 565876
rect 371844 565836 371850 565848
rect 373258 565836 373264 565848
rect 373316 565836 373322 565888
rect 516410 565836 516416 565888
rect 516468 565876 516474 565888
rect 521930 565876 521936 565888
rect 516468 565848 521936 565876
rect 516468 565836 516474 565848
rect 521930 565836 521936 565848
rect 521988 565836 521994 565888
rect 371786 564680 371792 564732
rect 371844 564720 371850 564732
rect 374270 564720 374276 564732
rect 371844 564692 374276 564720
rect 371844 564680 371850 564692
rect 374270 564680 374276 564692
rect 374328 564680 374334 564732
rect 516502 564680 516508 564732
rect 516560 564720 516566 564732
rect 520550 564720 520556 564732
rect 516560 564692 520556 564720
rect 516560 564680 516566 564692
rect 520550 564680 520556 564692
rect 520608 564680 520614 564732
rect 444374 564544 444380 564596
rect 444432 564584 444438 564596
rect 446490 564584 446496 564596
rect 444432 564556 446496 564584
rect 444432 564544 444438 564556
rect 446490 564544 446496 564556
rect 446548 564544 446554 564596
rect 516410 564476 516416 564528
rect 516468 564516 516474 564528
rect 519262 564516 519268 564528
rect 516468 564488 519268 564516
rect 516468 564476 516474 564488
rect 519262 564476 519268 564488
rect 519320 564476 519326 564528
rect 516318 563728 516324 563780
rect 516376 563768 516382 563780
rect 520274 563768 520280 563780
rect 516376 563740 520280 563768
rect 516376 563728 516382 563740
rect 520274 563728 520280 563740
rect 520332 563728 520338 563780
rect 516318 563252 516324 563304
rect 516376 563292 516382 563304
rect 518986 563292 518992 563304
rect 516376 563264 518992 563292
rect 516376 563252 516382 563264
rect 518986 563252 518992 563264
rect 519044 563252 519050 563304
rect 371786 563048 371792 563100
rect 371844 563088 371850 563100
rect 374362 563088 374368 563100
rect 371844 563060 374368 563088
rect 371844 563048 371850 563060
rect 374362 563048 374368 563060
rect 374420 563048 374426 563100
rect 445662 563048 445668 563100
rect 445720 563088 445726 563100
rect 450538 563088 450544 563100
rect 445720 563060 450544 563088
rect 445720 563048 445726 563060
rect 450538 563048 450544 563060
rect 450596 563048 450602 563100
rect 516318 563048 516324 563100
rect 516376 563088 516382 563100
rect 517790 563088 517796 563100
rect 516376 563060 517796 563088
rect 516376 563048 516382 563060
rect 517790 563048 517796 563060
rect 517848 563048 517854 563100
rect 371786 562504 371792 562556
rect 371844 562544 371850 562556
rect 374454 562544 374460 562556
rect 371844 562516 374460 562544
rect 371844 562504 371850 562516
rect 374454 562504 374460 562516
rect 374512 562504 374518 562556
rect 516318 562504 516324 562556
rect 516376 562544 516382 562556
rect 519078 562544 519084 562556
rect 516376 562516 519084 562544
rect 516376 562504 516382 562516
rect 519078 562504 519084 562516
rect 519136 562504 519142 562556
rect 516318 561960 516324 562012
rect 516376 562000 516382 562012
rect 517882 562000 517888 562012
rect 516376 561972 517888 562000
rect 516376 561960 516382 561972
rect 517882 561960 517888 561972
rect 517940 561960 517946 562012
rect 516318 561416 516324 561468
rect 516376 561456 516382 561468
rect 517974 561456 517980 561468
rect 516376 561428 517980 561456
rect 516376 561416 516382 561428
rect 517974 561416 517980 561428
rect 518032 561416 518038 561468
rect 444374 561144 444380 561196
rect 444432 561184 444438 561196
rect 446582 561184 446588 561196
rect 444432 561156 446588 561184
rect 444432 561144 444438 561156
rect 446582 561144 446588 561156
rect 446640 561144 446646 561196
rect 371786 560872 371792 560924
rect 371844 560912 371850 560924
rect 375558 560912 375564 560924
rect 371844 560884 375564 560912
rect 371844 560872 371850 560884
rect 375558 560872 375564 560884
rect 375616 560872 375622 560924
rect 371786 560328 371792 560380
rect 371844 560368 371850 560380
rect 376110 560368 376116 560380
rect 371844 560340 376116 560368
rect 371844 560328 371850 560340
rect 376110 560328 376116 560340
rect 376168 560328 376174 560380
rect 371786 559104 371792 559156
rect 371844 559144 371850 559156
rect 374546 559144 374552 559156
rect 371844 559116 374552 559144
rect 371844 559104 371850 559116
rect 374546 559104 374552 559116
rect 374604 559104 374610 559156
rect 516318 558968 516324 559020
rect 516376 559008 516382 559020
rect 524690 559008 524696 559020
rect 516376 558980 524696 559008
rect 516376 558968 516382 558980
rect 524690 558968 524696 558980
rect 524748 558968 524754 559020
rect 371878 558900 371884 558952
rect 371936 558940 371942 558952
rect 377122 558940 377128 558952
rect 371936 558912 377128 558940
rect 371936 558900 371942 558912
rect 377122 558900 377128 558912
rect 377180 558900 377186 558952
rect 516502 558900 516508 558952
rect 516560 558940 516566 558952
rect 525794 558940 525800 558952
rect 516560 558912 525800 558940
rect 516560 558900 516566 558912
rect 525794 558900 525800 558912
rect 525852 558900 525858 558952
rect 371786 558152 371792 558204
rect 371844 558192 371850 558204
rect 374086 558192 374092 558204
rect 371844 558164 374092 558192
rect 371844 558152 371850 558164
rect 374086 558152 374092 558164
rect 374144 558152 374150 558204
rect 371786 558016 371792 558068
rect 371844 558056 371850 558068
rect 375650 558056 375656 558068
rect 371844 558028 375656 558056
rect 371844 558016 371850 558028
rect 375650 558016 375656 558028
rect 375708 558056 375714 558068
rect 441614 558056 441620 558068
rect 375708 558028 441620 558056
rect 375708 558016 375714 558028
rect 441614 558016 441620 558028
rect 441672 558016 441678 558068
rect 516502 557744 516508 557796
rect 516560 557784 516566 557796
rect 519170 557784 519176 557796
rect 516560 557756 519176 557784
rect 516560 557744 516566 557756
rect 519170 557744 519176 557756
rect 519228 557744 519234 557796
rect 516318 557676 516324 557728
rect 516376 557716 516382 557728
rect 523034 557716 523040 557728
rect 516376 557688 523040 557716
rect 516376 557676 516382 557688
rect 523034 557676 523040 557688
rect 523092 557676 523098 557728
rect 444374 557608 444380 557660
rect 444432 557648 444438 557660
rect 447134 557648 447140 557660
rect 444432 557620 447140 557648
rect 444432 557608 444438 557620
rect 447134 557608 447140 557620
rect 447192 557608 447198 557660
rect 516778 557608 516784 557660
rect 516836 557608 516842 557660
rect 517054 557608 517060 557660
rect 517112 557648 517118 557660
rect 521838 557648 521844 557660
rect 517112 557620 521844 557648
rect 517112 557608 517118 557620
rect 521838 557608 521844 557620
rect 521896 557608 521902 557660
rect 516594 557540 516600 557592
rect 516652 557580 516658 557592
rect 516796 557580 516824 557608
rect 516652 557552 516824 557580
rect 516652 557540 516658 557552
rect 502978 557064 502984 557116
rect 503036 557104 503042 557116
rect 516134 557104 516140 557116
rect 503036 557076 516140 557104
rect 503036 557064 503042 557076
rect 516134 557064 516140 557076
rect 516192 557064 516198 557116
rect 501598 556996 501604 557048
rect 501656 557036 501662 557048
rect 516318 557036 516324 557048
rect 501656 557008 516324 557036
rect 501656 556996 501662 557008
rect 516318 556996 516324 557008
rect 516376 556996 516382 557048
rect 486418 556928 486424 556980
rect 486476 556968 486482 556980
rect 516594 556968 516600 556980
rect 486476 556940 516600 556968
rect 486476 556928 486482 556940
rect 516594 556928 516600 556940
rect 516652 556928 516658 556980
rect 454678 556860 454684 556912
rect 454736 556900 454742 556912
rect 516410 556900 516416 556912
rect 454736 556872 516416 556900
rect 454736 556860 454742 556872
rect 516410 556860 516416 556872
rect 516468 556860 516474 556912
rect 370498 556792 370504 556844
rect 370556 556832 370562 556844
rect 441706 556832 441712 556844
rect 370556 556804 441712 556832
rect 370556 556792 370562 556804
rect 441706 556792 441712 556804
rect 441764 556832 441770 556844
rect 513374 556832 513380 556844
rect 441764 556804 513380 556832
rect 441764 556792 441770 556804
rect 513374 556792 513380 556804
rect 513432 556792 513438 556844
rect 371786 556248 371792 556300
rect 371844 556288 371850 556300
rect 372890 556288 372896 556300
rect 371844 556260 372896 556288
rect 371844 556248 371850 556260
rect 372890 556248 372896 556260
rect 372948 556248 372954 556300
rect 516134 556248 516140 556300
rect 516192 556288 516198 556300
rect 521654 556288 521660 556300
rect 516192 556260 521660 556288
rect 516192 556248 516198 556260
rect 521654 556248 521660 556260
rect 521712 556248 521718 556300
rect 516226 556180 516232 556232
rect 516284 556220 516290 556232
rect 524506 556220 524512 556232
rect 516284 556192 524512 556220
rect 516284 556180 516290 556192
rect 524506 556180 524512 556192
rect 524564 556180 524570 556232
rect 376018 556112 376024 556164
rect 376076 556152 376082 556164
rect 516870 556152 516876 556164
rect 376076 556124 516876 556152
rect 376076 556112 376082 556124
rect 516870 556112 516876 556124
rect 516928 556112 516934 556164
rect 373258 556044 373264 556096
rect 373316 556084 373322 556096
rect 441614 556084 441620 556096
rect 373316 556056 441620 556084
rect 373316 556044 373322 556056
rect 441614 556044 441620 556056
rect 441672 556044 441678 556096
rect 376110 555976 376116 556028
rect 376168 556016 376174 556028
rect 444466 556016 444472 556028
rect 376168 555988 444472 556016
rect 376168 555976 376174 555988
rect 444466 555976 444472 555988
rect 444524 555976 444530 556028
rect 503346 555908 503352 555960
rect 503404 555948 503410 555960
rect 513466 555948 513472 555960
rect 503404 555920 513472 555948
rect 503404 555908 503410 555920
rect 513466 555908 513472 555920
rect 513524 555908 513530 555960
rect 503254 555840 503260 555892
rect 503312 555880 503318 555892
rect 513558 555880 513564 555892
rect 503312 555852 513564 555880
rect 503312 555840 503318 555852
rect 513558 555840 513564 555852
rect 513616 555840 513622 555892
rect 503162 555772 503168 555824
rect 503220 555812 503226 555824
rect 513650 555812 513656 555824
rect 503220 555784 513656 555812
rect 503220 555772 503226 555784
rect 513650 555772 513656 555784
rect 513708 555772 513714 555824
rect 503070 555704 503076 555756
rect 503128 555744 503134 555756
rect 513742 555744 513748 555756
rect 503128 555716 513748 555744
rect 503128 555704 503134 555716
rect 513742 555704 513748 555716
rect 513800 555704 513806 555756
rect 482278 555636 482284 555688
rect 482336 555676 482342 555688
rect 516502 555676 516508 555688
rect 482336 555648 516508 555676
rect 482336 555636 482342 555648
rect 516502 555636 516508 555648
rect 516560 555636 516566 555688
rect 464338 555568 464344 555620
rect 464396 555608 464402 555620
rect 516962 555608 516968 555620
rect 464396 555580 516968 555608
rect 464396 555568 464402 555580
rect 516962 555568 516968 555580
rect 517020 555568 517026 555620
rect 456702 555500 456708 555552
rect 456760 555540 456766 555552
rect 513834 555540 513840 555552
rect 456760 555512 513840 555540
rect 456760 555500 456766 555512
rect 513834 555500 513840 555512
rect 513892 555500 513898 555552
rect 449250 555432 449256 555484
rect 449308 555472 449314 555484
rect 516686 555472 516692 555484
rect 449308 555444 516692 555472
rect 449308 555432 449314 555444
rect 516686 555432 516692 555444
rect 516744 555432 516750 555484
rect 516778 554752 516784 554804
rect 516836 554792 516842 554804
rect 517514 554792 517520 554804
rect 516836 554764 517520 554792
rect 516836 554752 516842 554764
rect 517514 554752 517520 554764
rect 517572 554752 517578 554804
rect 435174 554684 435180 554736
rect 435232 554724 435238 554736
rect 506842 554724 506848 554736
rect 435232 554696 506848 554724
rect 435232 554684 435238 554696
rect 506842 554684 506848 554696
rect 506900 554684 506906 554736
rect 198642 554140 198648 554192
rect 198700 554180 198706 554192
rect 366910 554180 366916 554192
rect 198700 554152 366916 554180
rect 198700 554140 198706 554152
rect 366910 554140 366916 554152
rect 366968 554140 366974 554192
rect 302878 554072 302884 554124
rect 302936 554112 302942 554124
rect 510890 554112 510896 554124
rect 302936 554084 510896 554112
rect 302936 554072 302942 554084
rect 510890 554072 510896 554084
rect 510948 554072 510954 554124
rect 198550 554004 198556 554056
rect 198608 554044 198614 554056
rect 438946 554044 438952 554056
rect 198608 554016 438952 554044
rect 198608 554004 198614 554016
rect 438946 554004 438952 554016
rect 439004 554004 439010 554056
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 266446 553432 266452 553444
rect 3476 553404 266452 553432
rect 3476 553392 3482 553404
rect 266446 553392 266452 553404
rect 266504 553392 266510 553444
rect 512914 553392 512920 553444
rect 512972 553432 512978 553444
rect 514754 553432 514760 553444
rect 512972 553404 514760 553432
rect 512972 553392 512978 553404
rect 514754 553392 514760 553404
rect 514812 553392 514818 553444
rect 368934 551896 368940 551948
rect 368992 551936 368998 551948
rect 369302 551936 369308 551948
rect 368992 551908 369308 551936
rect 368992 551896 368998 551908
rect 369302 551896 369308 551908
rect 369360 551896 369366 551948
rect 448146 541628 448152 541680
rect 448204 541668 448210 541680
rect 521930 541668 521936 541680
rect 448204 541640 521936 541668
rect 448204 541628 448210 541640
rect 521930 541628 521936 541640
rect 521988 541628 521994 541680
rect 230382 536800 230388 536852
rect 230440 536840 230446 536852
rect 580166 536840 580172 536852
rect 230440 536812 580172 536840
rect 230440 536800 230446 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 448238 536052 448244 536104
rect 448296 536092 448302 536104
rect 520550 536092 520556 536104
rect 448296 536064 520556 536092
rect 448296 536052 448302 536064
rect 520550 536052 520556 536064
rect 520608 536052 520614 536104
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 267826 527184 267832 527196
rect 3476 527156 267832 527184
rect 3476 527144 3482 527156
rect 267826 527144 267832 527156
rect 267884 527144 267890 527196
rect 449158 526396 449164 526448
rect 449216 526436 449222 526448
rect 449342 526436 449348 526448
rect 449216 526408 449348 526436
rect 449216 526396 449222 526408
rect 449342 526396 449348 526408
rect 449400 526436 449406 526448
rect 517882 526436 517888 526448
rect 449400 526408 517888 526436
rect 449400 526396 449406 526408
rect 517882 526396 517888 526408
rect 517940 526396 517946 526448
rect 230290 524424 230296 524476
rect 230348 524464 230354 524476
rect 580166 524464 580172 524476
rect 230348 524436 580172 524464
rect 230348 524424 230354 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 446490 523676 446496 523728
rect 446548 523716 446554 523728
rect 525794 523716 525800 523728
rect 446548 523688 525800 523716
rect 446548 523676 446554 523688
rect 525794 523676 525800 523688
rect 525852 523676 525858 523728
rect 376202 522928 376208 522980
rect 376260 522968 376266 522980
rect 376662 522968 376668 522980
rect 376260 522940 376668 522968
rect 376260 522928 376266 522940
rect 376662 522928 376668 522940
rect 376720 522928 376726 522980
rect 450538 522316 450544 522368
rect 450596 522356 450602 522368
rect 524690 522356 524696 522368
rect 450596 522328 524696 522356
rect 450596 522316 450602 522328
rect 524690 522316 524696 522328
rect 524748 522316 524754 522368
rect 376662 522248 376668 522300
rect 376720 522288 376726 522300
rect 454034 522288 454040 522300
rect 376720 522260 454040 522288
rect 376720 522248 376726 522260
rect 454034 522248 454040 522260
rect 454092 522288 454098 522300
rect 454678 522288 454684 522300
rect 454092 522260 454684 522288
rect 454092 522248 454098 522260
rect 454678 522248 454684 522260
rect 454736 522248 454742 522300
rect 448054 520888 448060 520940
rect 448112 520928 448118 520940
rect 517790 520928 517796 520940
rect 448112 520900 517796 520928
rect 448112 520888 448118 520900
rect 517790 520888 517796 520900
rect 517848 520888 517854 520940
rect 447870 517828 447876 517880
rect 447928 517868 447934 517880
rect 448422 517868 448428 517880
rect 447928 517840 448428 517868
rect 447928 517828 447934 517840
rect 448422 517828 448428 517840
rect 448480 517828 448486 517880
rect 448422 517488 448428 517540
rect 448480 517528 448486 517540
rect 516410 517528 516416 517540
rect 448480 517500 516416 517528
rect 448480 517488 448486 517500
rect 516410 517488 516416 517500
rect 516468 517528 516474 517540
rect 520458 517528 520464 517540
rect 516468 517500 520464 517528
rect 516468 517488 516474 517500
rect 520458 517488 520464 517500
rect 520516 517488 520522 517540
rect 369118 516944 369124 516996
rect 369176 516984 369182 516996
rect 369486 516984 369492 516996
rect 369176 516956 369492 516984
rect 369176 516944 369182 516956
rect 369486 516944 369492 516956
rect 369544 516944 369550 516996
rect 516134 516060 516140 516112
rect 516192 516100 516198 516112
rect 519262 516100 519268 516112
rect 516192 516072 519268 516100
rect 516192 516060 516198 516072
rect 519262 516060 519268 516072
rect 519320 516060 519326 516112
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 270494 514808 270500 514820
rect 3476 514780 270500 514808
rect 3476 514768 3482 514780
rect 270494 514768 270500 514780
rect 270552 514768 270558 514820
rect 447870 514768 447876 514820
rect 447928 514808 447934 514820
rect 516134 514808 516140 514820
rect 447928 514780 516140 514808
rect 447928 514768 447934 514780
rect 516134 514768 516140 514780
rect 516192 514768 516198 514820
rect 507854 514020 507860 514072
rect 507912 514060 507918 514072
rect 513374 514060 513380 514072
rect 507912 514032 513380 514060
rect 507912 514020 507918 514032
rect 513374 514020 513380 514032
rect 513432 514020 513438 514072
rect 517146 514020 517152 514072
rect 517204 514060 517210 514072
rect 518158 514060 518164 514072
rect 517204 514032 518164 514060
rect 517204 514020 517210 514032
rect 518158 514020 518164 514032
rect 518216 514060 518222 514072
rect 524598 514060 524604 514072
rect 518216 514032 524604 514060
rect 518216 514020 518222 514032
rect 524598 514020 524604 514032
rect 524656 514020 524662 514072
rect 444374 513748 444380 513800
rect 444432 513788 444438 513800
rect 444926 513788 444932 513800
rect 444432 513760 444932 513788
rect 444432 513748 444438 513760
rect 444926 513748 444932 513760
rect 444984 513788 444990 513800
rect 446398 513788 446404 513800
rect 444984 513760 446404 513788
rect 444984 513748 444990 513760
rect 446398 513748 446404 513760
rect 446456 513748 446462 513800
rect 444558 512728 444564 512780
rect 444616 512768 444622 512780
rect 483658 512768 483664 512780
rect 444616 512740 483664 512768
rect 444616 512728 444622 512740
rect 483658 512728 483664 512740
rect 483716 512728 483722 512780
rect 516134 512728 516140 512780
rect 516192 512768 516198 512780
rect 520366 512768 520372 512780
rect 516192 512740 520372 512768
rect 516192 512728 516198 512740
rect 520366 512728 520372 512740
rect 520424 512728 520430 512780
rect 447778 512660 447784 512712
rect 447836 512700 447842 512712
rect 513742 512700 513748 512712
rect 447836 512672 513748 512700
rect 447836 512660 447842 512672
rect 513742 512660 513748 512672
rect 513800 512660 513806 512712
rect 445386 512592 445392 512644
rect 445444 512632 445450 512644
rect 514846 512632 514852 512644
rect 445444 512604 514852 512632
rect 445444 512592 445450 512604
rect 514846 512592 514852 512604
rect 514904 512592 514910 512644
rect 445662 511912 445668 511964
rect 445720 511952 445726 511964
rect 485038 511952 485044 511964
rect 445720 511924 485044 511952
rect 445720 511912 445726 511924
rect 485038 511912 485044 511924
rect 485096 511912 485102 511964
rect 369118 511776 369124 511828
rect 369176 511816 369182 511828
rect 369394 511816 369400 511828
rect 369176 511788 369400 511816
rect 369176 511776 369182 511788
rect 369394 511776 369400 511788
rect 369452 511776 369458 511828
rect 370958 511164 370964 511216
rect 371016 511204 371022 511216
rect 372982 511204 372988 511216
rect 371016 511176 372988 511204
rect 371016 511164 371022 511176
rect 372982 511164 372988 511176
rect 373040 511164 373046 511216
rect 517698 510620 517704 510672
rect 517756 510660 517762 510672
rect 518894 510660 518900 510672
rect 517756 510632 518900 510660
rect 517756 510620 517762 510632
rect 518894 510620 518900 510632
rect 518952 510620 518958 510672
rect 370958 510008 370964 510060
rect 371016 510048 371022 510060
rect 374638 510048 374644 510060
rect 371016 510020 374644 510048
rect 371016 510008 371022 510020
rect 374638 510008 374644 510020
rect 374696 510048 374702 510060
rect 374914 510048 374920 510060
rect 374696 510020 374920 510048
rect 374696 510008 374702 510020
rect 374914 510008 374920 510020
rect 374972 510008 374978 510060
rect 445662 509940 445668 509992
rect 445720 509980 445726 509992
rect 452654 509980 452660 509992
rect 445720 509952 452660 509980
rect 445720 509940 445726 509952
rect 452654 509940 452660 509952
rect 452712 509980 452718 509992
rect 489178 509980 489184 509992
rect 452712 509952 489184 509980
rect 452712 509940 452718 509952
rect 489178 509940 489184 509952
rect 489236 509940 489242 509992
rect 445570 509872 445576 509924
rect 445628 509912 445634 509924
rect 451274 509912 451280 509924
rect 445628 509884 451280 509912
rect 445628 509872 445634 509884
rect 451274 509872 451280 509884
rect 451332 509912 451338 509924
rect 490558 509912 490564 509924
rect 451332 509884 490564 509912
rect 451332 509872 451338 509884
rect 490558 509872 490564 509884
rect 490616 509872 490622 509924
rect 516134 509872 516140 509924
rect 516192 509912 516198 509924
rect 521746 509912 521752 509924
rect 516192 509884 521752 509912
rect 516192 509872 516198 509884
rect 521746 509872 521752 509884
rect 521804 509872 521810 509924
rect 516134 508784 516140 508836
rect 516192 508824 516198 508836
rect 519354 508824 519360 508836
rect 516192 508796 519360 508824
rect 516192 508784 516198 508796
rect 519354 508784 519360 508796
rect 519412 508784 519418 508836
rect 445662 508512 445668 508564
rect 445720 508552 445726 508564
rect 450170 508552 450176 508564
rect 445720 508524 450176 508552
rect 445720 508512 445726 508524
rect 450170 508512 450176 508524
rect 450228 508552 450234 508564
rect 493318 508552 493324 508564
rect 450228 508524 493324 508552
rect 450228 508512 450234 508524
rect 493318 508512 493324 508524
rect 493376 508512 493382 508564
rect 445570 507832 445576 507884
rect 445628 507872 445634 507884
rect 445628 507844 448560 507872
rect 445628 507832 445634 507844
rect 448532 507804 448560 507844
rect 519354 507832 519360 507884
rect 519412 507872 519418 507884
rect 520642 507872 520648 507884
rect 519412 507844 520648 507872
rect 519412 507832 519418 507844
rect 520642 507832 520648 507844
rect 520700 507832 520706 507884
rect 449158 507804 449164 507816
rect 448532 507776 449164 507804
rect 449158 507764 449164 507776
rect 449216 507804 449222 507816
rect 503346 507804 503352 507816
rect 449216 507776 503352 507804
rect 449216 507764 449222 507776
rect 503346 507764 503352 507776
rect 503404 507764 503410 507816
rect 516134 507764 516140 507816
rect 516192 507804 516198 507816
rect 521930 507804 521936 507816
rect 516192 507776 521936 507804
rect 516192 507764 516198 507776
rect 521930 507764 521936 507776
rect 521988 507764 521994 507816
rect 445570 507152 445576 507204
rect 445628 507192 445634 507204
rect 450078 507192 450084 507204
rect 445628 507164 450084 507192
rect 445628 507152 445634 507164
rect 450078 507152 450084 507164
rect 450136 507192 450142 507204
rect 497458 507192 497464 507204
rect 450136 507164 497464 507192
rect 450136 507152 450142 507164
rect 497458 507152 497464 507164
rect 497516 507152 497522 507204
rect 445662 507084 445668 507136
rect 445720 507124 445726 507136
rect 449986 507124 449992 507136
rect 445720 507096 449992 507124
rect 445720 507084 445726 507096
rect 449986 507084 449992 507096
rect 450044 507124 450050 507136
rect 500218 507124 500224 507136
rect 450044 507096 500224 507124
rect 450044 507084 450050 507096
rect 500218 507084 500224 507096
rect 500276 507084 500282 507136
rect 370958 506472 370964 506524
rect 371016 506512 371022 506524
rect 374178 506512 374184 506524
rect 371016 506484 374184 506512
rect 371016 506472 371022 506484
rect 374178 506472 374184 506484
rect 374236 506512 374242 506524
rect 374822 506512 374828 506524
rect 374236 506484 374828 506512
rect 374236 506472 374242 506484
rect 374822 506472 374828 506484
rect 374880 506472 374886 506524
rect 445570 505860 445576 505912
rect 445628 505900 445634 505912
rect 448514 505900 448520 505912
rect 445628 505872 448520 505900
rect 445628 505860 445634 505872
rect 448514 505860 448520 505872
rect 448572 505900 448578 505912
rect 449250 505900 449256 505912
rect 448572 505872 449256 505900
rect 448572 505860 448578 505872
rect 449250 505860 449256 505872
rect 449308 505860 449314 505912
rect 369118 505520 369124 505572
rect 369176 505560 369182 505572
rect 369486 505560 369492 505572
rect 369176 505532 369492 505560
rect 369176 505520 369182 505532
rect 369486 505520 369492 505532
rect 369544 505520 369550 505572
rect 370038 505452 370044 505504
rect 370096 505492 370102 505504
rect 373258 505492 373264 505504
rect 370096 505464 373264 505492
rect 370096 505452 370102 505464
rect 373258 505452 373264 505464
rect 373316 505452 373322 505504
rect 516962 505384 516968 505436
rect 517020 505424 517026 505436
rect 517606 505424 517612 505436
rect 517020 505396 517612 505424
rect 517020 505384 517026 505396
rect 517606 505384 517612 505396
rect 517664 505424 517670 505436
rect 520366 505424 520372 505436
rect 517664 505396 520372 505424
rect 517664 505384 517670 505396
rect 520366 505384 520372 505396
rect 520424 505384 520430 505436
rect 445662 505112 445668 505164
rect 445720 505152 445726 505164
rect 449894 505152 449900 505164
rect 445720 505124 449900 505152
rect 445720 505112 445726 505124
rect 449894 505112 449900 505124
rect 449952 505112 449958 505164
rect 448422 505044 448428 505096
rect 448480 505084 448486 505096
rect 452746 505084 452752 505096
rect 448480 505056 452752 505084
rect 448480 505044 448486 505056
rect 452746 505044 452752 505056
rect 452804 505044 452810 505096
rect 503254 505084 503260 505096
rect 460906 505056 503260 505084
rect 449894 504976 449900 505028
rect 449952 505016 449958 505028
rect 450538 505016 450544 505028
rect 449952 504988 450544 505016
rect 449952 504976 449958 504988
rect 450538 504976 450544 504988
rect 450596 505016 450602 505028
rect 460906 505016 460934 505056
rect 503254 505044 503260 505056
rect 503312 505044 503318 505096
rect 516134 505044 516140 505096
rect 516192 505084 516198 505096
rect 520550 505084 520556 505096
rect 516192 505056 520556 505084
rect 516192 505044 516198 505056
rect 520550 505044 520556 505056
rect 520608 505044 520614 505096
rect 450596 504988 460934 505016
rect 450596 504976 450602 504988
rect 458174 504432 458180 504484
rect 458232 504472 458238 504484
rect 464338 504472 464344 504484
rect 458232 504444 464344 504472
rect 458232 504432 458238 504444
rect 464338 504432 464344 504444
rect 464396 504432 464402 504484
rect 445662 504364 445668 504416
rect 445720 504404 445726 504416
rect 448606 504404 448612 504416
rect 445720 504376 448612 504404
rect 445720 504364 445726 504376
rect 448606 504364 448612 504376
rect 448664 504404 448670 504416
rect 501598 504404 501604 504416
rect 448664 504376 501604 504404
rect 448664 504364 448670 504376
rect 501598 504364 501604 504376
rect 501656 504364 501662 504416
rect 370958 504160 370964 504212
rect 371016 504200 371022 504212
rect 372614 504200 372620 504212
rect 371016 504172 372620 504200
rect 371016 504160 371022 504172
rect 372614 504160 372620 504172
rect 372672 504200 372678 504212
rect 373074 504200 373080 504212
rect 372672 504172 373080 504200
rect 372672 504160 372678 504172
rect 373074 504160 373080 504172
rect 373132 504160 373138 504212
rect 445294 503684 445300 503736
rect 445352 503724 445358 503736
rect 458174 503724 458180 503736
rect 445352 503696 458180 503724
rect 445352 503684 445358 503696
rect 458174 503684 458180 503696
rect 458232 503724 458238 503736
rect 458818 503724 458824 503736
rect 458232 503696 458824 503724
rect 458232 503684 458238 503696
rect 458818 503684 458824 503696
rect 458876 503684 458882 503736
rect 446398 503616 446404 503668
rect 446456 503656 446462 503668
rect 447870 503656 447876 503668
rect 446456 503628 447876 503656
rect 446456 503616 446462 503628
rect 447870 503616 447876 503628
rect 447928 503616 447934 503668
rect 370958 503140 370964 503192
rect 371016 503180 371022 503192
rect 374270 503180 374276 503192
rect 371016 503152 374276 503180
rect 371016 503140 371022 503152
rect 374270 503140 374276 503152
rect 374328 503140 374334 503192
rect 445202 502256 445208 502308
rect 445260 502296 445266 502308
rect 503162 502296 503168 502308
rect 445260 502268 503168 502296
rect 445260 502256 445266 502268
rect 503162 502256 503168 502268
rect 503220 502256 503226 502308
rect 459554 501576 459560 501628
rect 459612 501616 459618 501628
rect 460198 501616 460204 501628
rect 459612 501588 460204 501616
rect 459612 501576 459618 501588
rect 460198 501576 460204 501588
rect 460256 501616 460262 501628
rect 486418 501616 486424 501628
rect 460256 501588 486424 501616
rect 460256 501576 460262 501588
rect 486418 501576 486424 501588
rect 486476 501576 486482 501628
rect 516870 501372 516876 501424
rect 516928 501412 516934 501424
rect 518250 501412 518256 501424
rect 516928 501384 518256 501412
rect 516928 501372 516934 501384
rect 518250 501372 518256 501384
rect 518308 501412 518314 501424
rect 520274 501412 520280 501424
rect 518308 501384 520280 501412
rect 518308 501372 518314 501384
rect 520274 501372 520280 501384
rect 520332 501372 520338 501424
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 269114 501004 269120 501016
rect 3108 500976 269120 501004
rect 3108 500964 3114 500976
rect 269114 500964 269120 500976
rect 269172 500964 269178 501016
rect 445294 500964 445300 501016
rect 445352 501004 445358 501016
rect 459554 501004 459560 501016
rect 445352 500976 459560 501004
rect 445352 500964 445358 500976
rect 459554 500964 459560 500976
rect 459612 500964 459618 501016
rect 445478 500896 445484 500948
rect 445536 500936 445542 500948
rect 503070 500936 503076 500948
rect 445536 500908 503076 500936
rect 445536 500896 445542 500908
rect 503070 500896 503076 500908
rect 503128 500896 503134 500948
rect 445570 500828 445576 500880
rect 445628 500868 445634 500880
rect 482278 500868 482284 500880
rect 445628 500840 482284 500868
rect 445628 500828 445634 500840
rect 482278 500828 482284 500840
rect 482336 500828 482342 500880
rect 445662 500760 445668 500812
rect 445720 500800 445726 500812
rect 456702 500800 456708 500812
rect 445720 500772 456708 500800
rect 445720 500760 445726 500772
rect 456702 500760 456708 500772
rect 456760 500760 456766 500812
rect 516134 500760 516140 500812
rect 516192 500800 516198 500812
rect 518986 500800 518992 500812
rect 516192 500772 518992 500800
rect 516192 500760 516198 500772
rect 518986 500760 518992 500772
rect 519044 500760 519050 500812
rect 516134 500488 516140 500540
rect 516192 500528 516198 500540
rect 517790 500528 517796 500540
rect 516192 500500 517796 500528
rect 516192 500488 516198 500500
rect 517790 500488 517796 500500
rect 517848 500488 517854 500540
rect 456702 500352 456708 500404
rect 456760 500392 456766 500404
rect 457438 500392 457444 500404
rect 456760 500364 457444 500392
rect 456760 500352 456766 500364
rect 457438 500352 457444 500364
rect 457496 500352 457502 500404
rect 372706 500284 372712 500336
rect 372764 500324 372770 500336
rect 373258 500324 373264 500336
rect 372764 500296 373264 500324
rect 372764 500284 372770 500296
rect 373258 500284 373264 500296
rect 373316 500284 373322 500336
rect 370958 499604 370964 499656
rect 371016 499644 371022 499656
rect 374362 499644 374368 499656
rect 371016 499616 374368 499644
rect 371016 499604 371022 499616
rect 374362 499604 374368 499616
rect 374420 499604 374426 499656
rect 444650 499468 444656 499520
rect 444708 499508 444714 499520
rect 454034 499508 454040 499520
rect 444708 499480 454040 499508
rect 444708 499468 444714 499480
rect 454034 499468 454040 499480
rect 454092 499468 454098 499520
rect 466822 498788 466828 498840
rect 466880 498828 466886 498840
rect 467742 498828 467748 498840
rect 466880 498800 467748 498828
rect 466880 498788 466886 498800
rect 467742 498788 467748 498800
rect 467800 498828 467806 498840
rect 502978 498828 502984 498840
rect 467800 498800 502984 498828
rect 467800 498788 467806 498800
rect 502978 498788 502984 498800
rect 503036 498788 503042 498840
rect 370958 498448 370964 498500
rect 371016 498488 371022 498500
rect 374454 498488 374460 498500
rect 371016 498460 374460 498488
rect 371016 498448 371022 498460
rect 374454 498448 374460 498460
rect 374512 498448 374518 498500
rect 516134 498448 516140 498500
rect 516192 498488 516198 498500
rect 519078 498488 519084 498500
rect 516192 498460 519084 498488
rect 516192 498448 516198 498460
rect 519078 498448 519084 498460
rect 519136 498448 519142 498500
rect 445570 498176 445576 498228
rect 445628 498216 445634 498228
rect 466822 498216 466828 498228
rect 445628 498188 466828 498216
rect 445628 498176 445634 498188
rect 466822 498176 466828 498188
rect 466880 498176 466886 498228
rect 516134 498108 516140 498160
rect 516192 498148 516198 498160
rect 517882 498148 517888 498160
rect 516192 498120 517888 498148
rect 516192 498108 516198 498120
rect 517882 498108 517888 498120
rect 517940 498108 517946 498160
rect 445478 497768 445484 497820
rect 445536 497808 445542 497820
rect 449250 497808 449256 497820
rect 445536 497780 449256 497808
rect 445536 497768 445542 497780
rect 449250 497768 449256 497780
rect 449308 497768 449314 497820
rect 445570 496952 445576 497004
rect 445628 496992 445634 497004
rect 447502 496992 447508 497004
rect 445628 496964 447508 496992
rect 445628 496952 445634 496964
rect 447502 496952 447508 496964
rect 447560 496952 447566 497004
rect 445754 496816 445760 496868
rect 445812 496856 445818 496868
rect 446306 496856 446312 496868
rect 445812 496828 446312 496856
rect 445812 496816 445818 496828
rect 446306 496816 446312 496828
rect 446364 496816 446370 496868
rect 447134 496816 447140 496868
rect 447192 496856 447198 496868
rect 449342 496856 449348 496868
rect 447192 496828 449348 496856
rect 447192 496816 447198 496828
rect 449342 496816 449348 496828
rect 449400 496816 449406 496868
rect 516226 495456 516232 495508
rect 516284 495496 516290 495508
rect 517514 495496 517520 495508
rect 516284 495468 517520 495496
rect 516284 495456 516290 495468
rect 517514 495456 517520 495468
rect 517572 495496 517578 495508
rect 517974 495496 517980 495508
rect 517572 495468 517980 495496
rect 517572 495456 517578 495468
rect 517974 495456 517980 495468
rect 518032 495456 518038 495508
rect 370958 494776 370964 494828
rect 371016 494816 371022 494828
rect 375558 494816 375564 494828
rect 371016 494788 375564 494816
rect 371016 494776 371022 494788
rect 375558 494776 375564 494788
rect 375616 494816 375622 494828
rect 376202 494816 376208 494828
rect 375616 494788 376208 494816
rect 375616 494776 375622 494788
rect 376202 494776 376208 494788
rect 376260 494776 376266 494828
rect 445294 494708 445300 494760
rect 445352 494748 445358 494760
rect 445570 494748 445576 494760
rect 445352 494720 445576 494748
rect 445352 494708 445358 494720
rect 445570 494708 445576 494720
rect 445628 494708 445634 494760
rect 445294 494572 445300 494624
rect 445352 494612 445358 494624
rect 446122 494612 446128 494624
rect 445352 494584 446128 494612
rect 445352 494572 445358 494584
rect 446122 494572 446128 494584
rect 446180 494612 446186 494624
rect 448146 494612 448152 494624
rect 446180 494584 448152 494612
rect 446180 494572 446186 494584
rect 448146 494572 448152 494584
rect 448204 494572 448210 494624
rect 442442 494028 442448 494080
rect 442500 494068 442506 494080
rect 442902 494068 442908 494080
rect 442500 494040 442908 494068
rect 442500 494028 442506 494040
rect 442902 494028 442908 494040
rect 442960 494068 442966 494080
rect 452746 494068 452752 494080
rect 442960 494040 452752 494068
rect 442960 494028 442966 494040
rect 452746 494028 452752 494040
rect 452804 494028 452810 494080
rect 370958 493960 370964 494012
rect 371016 494000 371022 494012
rect 375558 494000 375564 494012
rect 371016 493972 375564 494000
rect 371016 493960 371022 493972
rect 375558 493960 375564 493972
rect 375616 494000 375622 494012
rect 376110 494000 376116 494012
rect 375616 493972 376116 494000
rect 375616 493960 375622 493972
rect 376110 493960 376116 493972
rect 376168 493960 376174 494012
rect 446214 493960 446220 494012
rect 446272 494000 446278 494012
rect 448238 494000 448244 494012
rect 446272 493972 448244 494000
rect 446272 493960 446278 493972
rect 448238 493960 448244 493972
rect 448296 493960 448302 494012
rect 516226 493960 516232 494012
rect 516284 494000 516290 494012
rect 525794 494000 525800 494012
rect 516284 493972 525800 494000
rect 516284 493960 516290 493972
rect 525794 493960 525800 493972
rect 525852 493960 525858 494012
rect 445294 493348 445300 493400
rect 445352 493388 445358 493400
rect 446214 493388 446220 493400
rect 445352 493360 446220 493388
rect 445352 493348 445358 493360
rect 446214 493348 446220 493360
rect 446272 493348 446278 493400
rect 370774 493280 370780 493332
rect 370832 493320 370838 493332
rect 377122 493320 377128 493332
rect 370832 493292 377128 493320
rect 370832 493280 370838 493292
rect 377122 493280 377128 493292
rect 377180 493280 377186 493332
rect 444650 493280 444656 493332
rect 444708 493320 444714 493332
rect 446398 493320 446404 493332
rect 444708 493292 446404 493320
rect 444708 493280 444714 493292
rect 446398 493280 446404 493292
rect 446456 493320 446462 493332
rect 446950 493320 446956 493332
rect 446456 493292 446956 493320
rect 446456 493280 446462 493292
rect 446950 493280 446956 493292
rect 447008 493280 447014 493332
rect 516134 492600 516140 492652
rect 516192 492640 516198 492652
rect 524690 492640 524696 492652
rect 516192 492612 524696 492640
rect 516192 492600 516198 492612
rect 524690 492600 524696 492612
rect 524748 492600 524754 492652
rect 370866 492328 370872 492380
rect 370924 492368 370930 492380
rect 374546 492368 374552 492380
rect 370924 492340 374552 492368
rect 370924 492328 370930 492340
rect 374546 492328 374552 492340
rect 374604 492368 374610 492380
rect 377214 492368 377220 492380
rect 374604 492340 377220 492368
rect 374604 492328 374610 492340
rect 377214 492328 377220 492340
rect 377272 492328 377278 492380
rect 448790 491648 448796 491700
rect 448848 491688 448854 491700
rect 450630 491688 450636 491700
rect 448848 491660 450636 491688
rect 448848 491648 448854 491660
rect 450630 491648 450636 491660
rect 450688 491648 450694 491700
rect 369118 491308 369124 491360
rect 369176 491348 369182 491360
rect 369302 491348 369308 491360
rect 369176 491320 369308 491348
rect 369176 491308 369182 491320
rect 369302 491308 369308 491320
rect 369360 491308 369366 491360
rect 443546 491308 443552 491360
rect 443604 491348 443610 491360
rect 443604 491320 444420 491348
rect 443604 491308 443610 491320
rect 444392 491280 444420 491320
rect 445938 491280 445944 491292
rect 444392 491252 445944 491280
rect 445938 491240 445944 491252
rect 445996 491240 446002 491292
rect 443914 491172 443920 491224
rect 443972 491212 443978 491224
rect 447134 491212 447140 491224
rect 443972 491184 447140 491212
rect 443972 491172 443978 491184
rect 447134 491172 447140 491184
rect 447192 491172 447198 491224
rect 516134 491172 516140 491224
rect 516192 491212 516198 491224
rect 519170 491212 519176 491224
rect 516192 491184 519176 491212
rect 516192 491172 516198 491184
rect 519170 491172 519176 491184
rect 519228 491212 519234 491224
rect 522114 491212 522120 491224
rect 519228 491184 522120 491212
rect 519228 491172 519234 491184
rect 522114 491172 522120 491184
rect 522172 491172 522178 491224
rect 445294 491036 445300 491088
rect 445352 491076 445358 491088
rect 445938 491076 445944 491088
rect 445352 491048 445944 491076
rect 445352 491036 445358 491048
rect 445938 491036 445944 491048
rect 445996 491076 446002 491088
rect 448054 491076 448060 491088
rect 445996 491048 448060 491076
rect 445996 491036 446002 491048
rect 448054 491036 448060 491048
rect 448112 491036 448118 491088
rect 370958 490288 370964 490340
rect 371016 490328 371022 490340
rect 374086 490328 374092 490340
rect 371016 490300 374092 490328
rect 371016 490288 371022 490300
rect 374086 490288 374092 490300
rect 374144 490328 374150 490340
rect 374546 490328 374552 490340
rect 374144 490300 374552 490328
rect 374144 490288 374150 490300
rect 374546 490288 374552 490300
rect 374604 490288 374610 490340
rect 516686 489812 516692 489864
rect 516744 489852 516750 489864
rect 521838 489852 521844 489864
rect 516744 489824 521844 489852
rect 516744 489812 516750 489824
rect 521838 489812 521844 489824
rect 521896 489812 521902 489864
rect 370406 489336 370412 489388
rect 370464 489376 370470 489388
rect 370682 489376 370688 489388
rect 370464 489348 370688 489376
rect 370464 489336 370470 489348
rect 370682 489336 370688 489348
rect 370740 489336 370746 489388
rect 443086 488724 443092 488776
rect 443144 488764 443150 488776
rect 447410 488764 447416 488776
rect 443144 488736 447416 488764
rect 443144 488724 443150 488736
rect 447410 488724 447416 488736
rect 447468 488724 447474 488776
rect 441890 488520 441896 488572
rect 441948 488560 441954 488572
rect 442350 488560 442356 488572
rect 441948 488532 442356 488560
rect 441948 488520 441954 488532
rect 442350 488520 442356 488532
rect 442408 488520 442414 488572
rect 517238 488452 517244 488504
rect 517296 488492 517302 488504
rect 523034 488492 523040 488504
rect 517296 488464 523040 488492
rect 517296 488452 517302 488464
rect 523034 488452 523040 488464
rect 523092 488452 523098 488504
rect 369394 488044 369400 488096
rect 369452 488084 369458 488096
rect 369762 488084 369768 488096
rect 369452 488056 369768 488084
rect 369452 488044 369458 488056
rect 369762 488044 369768 488056
rect 369820 488084 369826 488096
rect 375650 488084 375656 488096
rect 369820 488056 375656 488084
rect 369820 488044 369826 488056
rect 375650 488044 375656 488056
rect 375708 488044 375714 488096
rect 444650 487840 444656 487892
rect 444708 487880 444714 487892
rect 446490 487880 446496 487892
rect 444708 487852 446496 487880
rect 444708 487840 444714 487852
rect 446490 487840 446496 487852
rect 446548 487840 446554 487892
rect 445294 487296 445300 487348
rect 445352 487336 445358 487348
rect 448790 487336 448796 487348
rect 445352 487308 448796 487336
rect 445352 487296 445358 487308
rect 448790 487296 448796 487308
rect 448848 487296 448854 487348
rect 445478 487160 445484 487212
rect 445536 487200 445542 487212
rect 448698 487200 448704 487212
rect 445536 487172 448704 487200
rect 445536 487160 445542 487172
rect 448698 487160 448704 487172
rect 448756 487160 448762 487212
rect 516134 486412 516140 486464
rect 516192 486452 516198 486464
rect 520918 486452 520924 486464
rect 516192 486424 520924 486452
rect 516192 486412 516198 486424
rect 520918 486412 520924 486424
rect 520976 486452 520982 486464
rect 524506 486452 524512 486464
rect 520976 486424 524512 486452
rect 520976 486412 520982 486424
rect 524506 486412 524512 486424
rect 524564 486412 524570 486464
rect 446582 486004 446588 486056
rect 446640 486044 446646 486056
rect 513466 486044 513472 486056
rect 446640 486016 513472 486044
rect 446640 486004 446646 486016
rect 513466 486004 513472 486016
rect 513524 486004 513530 486056
rect 445478 485800 445484 485852
rect 445536 485840 445542 485852
rect 445846 485840 445852 485852
rect 445536 485812 445852 485840
rect 445536 485800 445542 485812
rect 445846 485800 445852 485812
rect 445904 485840 445910 485852
rect 446582 485840 446588 485852
rect 445904 485812 446588 485840
rect 445904 485800 445910 485812
rect 446582 485800 446588 485812
rect 446640 485800 446646 485852
rect 445110 485732 445116 485784
rect 445168 485772 445174 485784
rect 513374 485772 513380 485784
rect 445168 485744 513380 485772
rect 445168 485732 445174 485744
rect 513374 485732 513380 485744
rect 513432 485732 513438 485784
rect 516134 485732 516140 485784
rect 516192 485772 516198 485784
rect 521654 485772 521660 485784
rect 516192 485744 521660 485772
rect 516192 485732 516198 485744
rect 521654 485732 521660 485744
rect 521712 485732 521718 485784
rect 370958 485256 370964 485308
rect 371016 485296 371022 485308
rect 372890 485296 372896 485308
rect 371016 485268 372896 485296
rect 371016 485256 371022 485268
rect 372890 485256 372896 485268
rect 372948 485256 372954 485308
rect 447318 485052 447324 485104
rect 447376 485092 447382 485104
rect 513742 485092 513748 485104
rect 447376 485064 513748 485092
rect 447376 485052 447382 485064
rect 513742 485052 513748 485064
rect 513800 485052 513806 485104
rect 369118 484848 369124 484900
rect 369176 484848 369182 484900
rect 369136 484696 369164 484848
rect 369118 484644 369124 484696
rect 369176 484644 369182 484696
rect 445478 484576 445484 484628
rect 445536 484616 445542 484628
rect 447318 484616 447324 484628
rect 445536 484588 447324 484616
rect 445536 484576 445542 484588
rect 447318 484576 447324 484588
rect 447376 484576 447382 484628
rect 448698 484304 448704 484356
rect 448756 484344 448762 484356
rect 449342 484344 449348 484356
rect 448756 484316 449348 484344
rect 448756 484304 448762 484316
rect 449342 484304 449348 484316
rect 449400 484344 449406 484356
rect 516226 484344 516232 484356
rect 449400 484316 516232 484344
rect 449400 484304 449406 484316
rect 516226 484304 516232 484316
rect 516284 484304 516290 484356
rect 513098 484236 513104 484288
rect 513156 484276 513162 484288
rect 514754 484276 514760 484288
rect 513156 484248 514760 484276
rect 513156 484236 513162 484248
rect 514754 484236 514760 484248
rect 514812 484236 514818 484288
rect 444650 484168 444656 484220
rect 444708 484208 444714 484220
rect 447686 484208 447692 484220
rect 444708 484180 447692 484208
rect 444708 484168 444714 484180
rect 447686 484168 447692 484180
rect 447744 484168 447750 484220
rect 362862 482944 362868 482996
rect 362920 482984 362926 482996
rect 435174 482984 435180 482996
rect 362920 482956 435180 482984
rect 362920 482944 362926 482956
rect 435174 482944 435180 482956
rect 435232 482984 435238 482996
rect 506842 482984 506848 482996
rect 435232 482956 506848 482984
rect 435232 482944 435238 482956
rect 506842 482944 506848 482956
rect 506900 482944 506906 482996
rect 371142 482876 371148 482928
rect 371200 482916 371206 482928
rect 436738 482916 436744 482928
rect 371200 482888 436744 482916
rect 371200 482876 371206 482888
rect 436738 482876 436744 482888
rect 436796 482916 436802 482928
rect 508866 482916 508872 482928
rect 436796 482888 508872 482916
rect 436796 482876 436802 482888
rect 508866 482876 508872 482888
rect 508924 482916 508930 482928
rect 513558 482916 513564 482928
rect 508924 482888 513564 482916
rect 508924 482876 508930 482888
rect 513558 482876 513564 482888
rect 513616 482876 513622 482928
rect 369210 482808 369216 482860
rect 369268 482848 369274 482860
rect 369762 482848 369768 482860
rect 369268 482820 369768 482848
rect 369268 482808 369274 482820
rect 369762 482808 369768 482820
rect 369820 482848 369826 482860
rect 440970 482848 440976 482860
rect 369820 482820 440976 482848
rect 369820 482808 369826 482820
rect 440970 482808 440976 482820
rect 441028 482848 441034 482860
rect 512914 482848 512920 482860
rect 441028 482820 512920 482848
rect 441028 482808 441034 482820
rect 512914 482808 512920 482820
rect 512972 482808 512978 482860
rect 360838 482740 360844 482792
rect 360896 482780 360902 482792
rect 432966 482780 432972 482792
rect 360896 482752 432972 482780
rect 360896 482740 360902 482752
rect 432966 482740 432972 482752
rect 433024 482780 433030 482792
rect 504910 482780 504916 482792
rect 433024 482752 504916 482780
rect 433024 482740 433030 482752
rect 504910 482740 504916 482752
rect 504968 482740 504974 482792
rect 323578 482400 323584 482452
rect 323636 482440 323642 482452
rect 366910 482440 366916 482452
rect 323636 482412 366916 482440
rect 323636 482400 323642 482412
rect 366910 482400 366916 482412
rect 366968 482400 366974 482452
rect 302970 482332 302976 482384
rect 303028 482372 303034 482384
rect 438946 482372 438952 482384
rect 303028 482344 438952 482372
rect 303028 482332 303034 482344
rect 438946 482332 438952 482344
rect 439004 482332 439010 482384
rect 198458 482264 198464 482316
rect 198516 482304 198522 482316
rect 510890 482304 510896 482316
rect 198516 482276 510896 482304
rect 198516 482264 198522 482276
rect 510890 482264 510896 482276
rect 510948 482264 510954 482316
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 270586 474756 270592 474768
rect 3476 474728 270592 474756
rect 3476 474716 3482 474728
rect 270586 474716 270592 474728
rect 270644 474716 270650 474768
rect 227622 470568 227628 470620
rect 227680 470608 227686 470620
rect 580166 470608 580172 470620
rect 227680 470580 580172 470608
rect 227680 470568 227686 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 273254 462380 273260 462392
rect 3292 462352 273260 462380
rect 3292 462340 3298 462352
rect 273254 462340 273260 462352
rect 273312 462340 273318 462392
rect 445018 460164 445024 460216
rect 445076 460204 445082 460216
rect 516410 460204 516416 460216
rect 445076 460176 516416 460204
rect 445076 460164 445082 460176
rect 516410 460164 516416 460176
rect 516468 460164 516474 460216
rect 226150 456764 226156 456816
rect 226208 456804 226214 456816
rect 580166 456804 580172 456816
rect 226208 456776 580172 456804
rect 226208 456764 226214 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 373258 455404 373264 455456
rect 373316 455444 373322 455456
rect 373902 455444 373908 455456
rect 373316 455416 373908 455444
rect 373316 455404 373322 455416
rect 373902 455404 373908 455416
rect 373960 455444 373966 455456
rect 442074 455444 442080 455456
rect 373960 455416 442080 455444
rect 373960 455404 373966 455416
rect 442074 455404 442080 455416
rect 442132 455444 442138 455456
rect 443546 455444 443552 455456
rect 442132 455416 443552 455444
rect 442132 455404 442138 455416
rect 443546 455404 443552 455416
rect 443604 455404 443610 455456
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 271874 448576 271880 448588
rect 3200 448548 271880 448576
rect 3200 448536 3206 448548
rect 271874 448536 271880 448548
rect 271932 448536 271938 448588
rect 376202 447108 376208 447160
rect 376260 447148 376266 447160
rect 377306 447148 377312 447160
rect 376260 447120 377312 447148
rect 376260 447108 376266 447120
rect 377306 447108 377312 447120
rect 377364 447148 377370 447160
rect 442258 447148 442264 447160
rect 377364 447120 442264 447148
rect 377364 447108 377370 447120
rect 442258 447108 442264 447120
rect 442316 447148 442322 447160
rect 443454 447148 443460 447160
rect 442316 447120 443460 447148
rect 442316 447108 442322 447120
rect 443454 447108 443460 447120
rect 443512 447108 443518 447160
rect 445294 442892 445300 442944
rect 445352 442932 445358 442944
rect 445570 442932 445576 442944
rect 445352 442904 445576 442932
rect 445352 442892 445358 442904
rect 445570 442892 445576 442904
rect 445628 442892 445634 442944
rect 467098 442892 467104 442944
rect 467156 442932 467162 442944
rect 467742 442932 467748 442944
rect 467156 442904 467748 442932
rect 467156 442892 467162 442904
rect 467742 442892 467748 442904
rect 467800 442892 467806 442944
rect 376110 442280 376116 442332
rect 376168 442320 376174 442332
rect 376662 442320 376668 442332
rect 376168 442292 376668 442320
rect 376168 442280 376174 442292
rect 376662 442280 376668 442292
rect 376720 442280 376726 442332
rect 377490 442280 377496 442332
rect 377548 442320 377554 442332
rect 458818 442320 458824 442332
rect 377548 442292 458824 442320
rect 377548 442280 377554 442292
rect 458818 442280 458824 442292
rect 458876 442320 458882 442332
rect 513466 442320 513472 442332
rect 458876 442292 513472 442320
rect 458876 442280 458882 442292
rect 513466 442280 513472 442292
rect 513524 442280 513530 442332
rect 372062 442212 372068 442264
rect 372120 442252 372126 442264
rect 460198 442252 460204 442264
rect 372120 442224 460204 442252
rect 372120 442212 372126 442224
rect 460198 442212 460204 442224
rect 460256 442252 460262 442264
rect 516594 442252 516600 442264
rect 460256 442224 516600 442252
rect 460256 442212 460262 442224
rect 516594 442212 516600 442224
rect 516652 442212 516658 442264
rect 467098 441872 467104 441924
rect 467156 441912 467162 441924
rect 516686 441912 516692 441924
rect 467156 441884 516692 441912
rect 467156 441872 467162 441884
rect 516686 441872 516692 441884
rect 516744 441872 516750 441924
rect 457438 441804 457444 441856
rect 457496 441844 457502 441856
rect 516962 441844 516968 441856
rect 457496 441816 516968 441844
rect 457496 441804 457502 441816
rect 516962 441804 516968 441816
rect 517020 441804 517026 441856
rect 445294 441736 445300 441788
rect 445352 441776 445358 441788
rect 513374 441776 513380 441788
rect 445352 441748 513380 441776
rect 445352 441736 445358 441748
rect 513374 441736 513380 441748
rect 513432 441736 513438 441788
rect 445202 441668 445208 441720
rect 445260 441708 445266 441720
rect 516502 441708 516508 441720
rect 445260 441680 516508 441708
rect 445260 441668 445266 441680
rect 516502 441668 516508 441680
rect 516560 441668 516566 441720
rect 376110 441600 376116 441652
rect 376168 441640 376174 441652
rect 516226 441640 516232 441652
rect 376168 441612 516232 441640
rect 376168 441600 376174 441612
rect 516226 441600 516232 441612
rect 516284 441600 516290 441652
rect 516134 441532 516140 441584
rect 516192 441572 516198 441584
rect 524414 441572 524420 441584
rect 516192 441544 524420 441572
rect 516192 441532 516198 441544
rect 524414 441532 524420 441544
rect 524472 441532 524478 441584
rect 445110 441328 445116 441380
rect 445168 441368 445174 441380
rect 446306 441368 446312 441380
rect 445168 441340 446312 441368
rect 445168 441328 445174 441340
rect 446306 441328 446312 441340
rect 446364 441328 446370 441380
rect 446306 440376 446312 440428
rect 446364 440416 446370 440428
rect 447870 440416 447876 440428
rect 446364 440388 447876 440416
rect 446364 440376 446370 440388
rect 447870 440376 447876 440388
rect 447928 440376 447934 440428
rect 444466 440308 444472 440360
rect 444524 440348 444530 440360
rect 444524 440320 451274 440348
rect 444524 440308 444530 440320
rect 371234 440240 371240 440292
rect 371292 440280 371298 440292
rect 371418 440280 371424 440292
rect 371292 440252 371424 440280
rect 371292 440240 371298 440252
rect 371418 440240 371424 440252
rect 371476 440240 371482 440292
rect 445570 440240 445576 440292
rect 445628 440280 445634 440292
rect 447502 440280 447508 440292
rect 445628 440252 447508 440280
rect 445628 440240 445634 440252
rect 447502 440240 447508 440252
rect 447560 440280 447566 440292
rect 447778 440280 447784 440292
rect 447560 440252 447784 440280
rect 447560 440240 447566 440252
rect 447778 440240 447784 440252
rect 447836 440240 447842 440292
rect 451246 440280 451274 440320
rect 513742 440280 513748 440292
rect 451246 440252 513748 440280
rect 513742 440240 513748 440252
rect 513800 440240 513806 440292
rect 516870 439084 516876 439136
rect 516928 439124 516934 439136
rect 517698 439124 517704 439136
rect 516928 439096 517704 439124
rect 516928 439084 516934 439096
rect 517698 439084 517704 439096
rect 517756 439084 517762 439136
rect 444190 439016 444196 439068
rect 444248 439056 444254 439068
rect 447134 439056 447140 439068
rect 444248 439028 447140 439056
rect 444248 439016 444254 439028
rect 447134 439016 447140 439028
rect 447192 439016 447198 439068
rect 371786 438880 371792 438932
rect 371844 438920 371850 438932
rect 372154 438920 372160 438932
rect 371844 438892 372160 438920
rect 371844 438880 371850 438892
rect 372154 438880 372160 438892
rect 372212 438920 372218 438932
rect 378870 438920 378876 438932
rect 372212 438892 378876 438920
rect 372212 438880 372218 438892
rect 378870 438880 378876 438892
rect 378928 438880 378934 438932
rect 516134 438880 516140 438932
rect 516192 438920 516198 438932
rect 529934 438920 529940 438932
rect 516192 438892 529940 438920
rect 516192 438880 516198 438892
rect 529934 438880 529940 438892
rect 529992 438880 529998 438932
rect 371602 438132 371608 438184
rect 371660 438172 371666 438184
rect 378226 438172 378232 438184
rect 371660 438144 378232 438172
rect 371660 438132 371666 438144
rect 378226 438132 378232 438144
rect 378284 438132 378290 438184
rect 444650 437928 444656 437980
rect 444708 437968 444714 437980
rect 446030 437968 446036 437980
rect 444708 437940 446036 437968
rect 444708 437928 444714 437940
rect 446030 437928 446036 437940
rect 446088 437928 446094 437980
rect 516226 437520 516232 437572
rect 516284 437560 516290 437572
rect 524414 437560 524420 437572
rect 516284 437532 524420 437560
rect 516284 437520 516290 437532
rect 524414 437520 524420 437532
rect 524472 437520 524478 437572
rect 378226 437452 378232 437504
rect 378284 437492 378290 437504
rect 378962 437492 378968 437504
rect 378284 437464 378968 437492
rect 378284 437452 378290 437464
rect 378962 437452 378968 437464
rect 379020 437452 379026 437504
rect 380158 437492 380164 437504
rect 379900 437464 380164 437492
rect 371694 437384 371700 437436
rect 371752 437424 371758 437436
rect 372154 437424 372160 437436
rect 371752 437396 372160 437424
rect 371752 437384 371758 437396
rect 372154 437384 372160 437396
rect 372212 437384 372218 437436
rect 371786 437316 371792 437368
rect 371844 437356 371850 437368
rect 377030 437356 377036 437368
rect 371844 437328 377036 437356
rect 371844 437316 371850 437328
rect 377030 437316 377036 437328
rect 377088 437356 377094 437368
rect 378042 437356 378048 437368
rect 377088 437328 378048 437356
rect 377088 437316 377094 437328
rect 378042 437316 378048 437328
rect 378100 437316 378106 437368
rect 371602 437248 371608 437300
rect 371660 437288 371666 437300
rect 379900 437288 379928 437464
rect 380158 437452 380164 437464
rect 380216 437492 380222 437504
rect 399478 437492 399484 437504
rect 380216 437464 399484 437492
rect 380216 437452 380222 437464
rect 399478 437452 399484 437464
rect 399536 437452 399542 437504
rect 443638 437452 443644 437504
rect 443696 437492 443702 437504
rect 444374 437492 444380 437504
rect 443696 437464 444380 437492
rect 443696 437452 443702 437464
rect 444374 437452 444380 437464
rect 444432 437452 444438 437504
rect 446030 437452 446036 437504
rect 446088 437492 446094 437504
rect 446674 437492 446680 437504
rect 446088 437464 446680 437492
rect 446088 437452 446094 437464
rect 446674 437452 446680 437464
rect 446732 437452 446738 437504
rect 516134 437452 516140 437504
rect 516192 437492 516198 437504
rect 528738 437492 528744 437504
rect 516192 437464 528744 437492
rect 516192 437452 516198 437464
rect 528738 437452 528744 437464
rect 528796 437452 528802 437504
rect 371660 437260 379928 437288
rect 371660 437248 371666 437260
rect 516502 436840 516508 436892
rect 516560 436880 516566 436892
rect 516870 436880 516876 436892
rect 516560 436852 516876 436880
rect 516560 436840 516566 436852
rect 516870 436840 516876 436852
rect 516928 436840 516934 436892
rect 371694 436772 371700 436824
rect 371752 436812 371758 436824
rect 373994 436812 374000 436824
rect 371752 436784 374000 436812
rect 371752 436772 371758 436784
rect 373994 436772 374000 436784
rect 374052 436812 374058 436824
rect 379238 436812 379244 436824
rect 374052 436784 379244 436812
rect 374052 436772 374058 436784
rect 379238 436772 379244 436784
rect 379296 436772 379302 436824
rect 445110 436772 445116 436824
rect 445168 436812 445174 436824
rect 445294 436812 445300 436824
rect 445168 436784 445300 436812
rect 445168 436772 445174 436784
rect 445294 436772 445300 436784
rect 445352 436772 445358 436824
rect 378042 436704 378048 436756
rect 378100 436744 378106 436756
rect 387058 436744 387064 436756
rect 378100 436716 387064 436744
rect 378100 436704 378106 436716
rect 387058 436704 387064 436716
rect 387116 436704 387122 436756
rect 444374 436704 444380 436756
rect 444432 436744 444438 436756
rect 446582 436744 446588 436756
rect 444432 436716 446588 436744
rect 444432 436704 444438 436716
rect 446582 436704 446588 436716
rect 446640 436704 446646 436756
rect 516226 436228 516232 436280
rect 516284 436268 516290 436280
rect 523034 436268 523040 436280
rect 516284 436240 523040 436268
rect 516284 436228 516290 436240
rect 523034 436228 523040 436240
rect 523092 436228 523098 436280
rect 516502 436160 516508 436212
rect 516560 436200 516566 436212
rect 525794 436200 525800 436212
rect 516560 436172 525800 436200
rect 516560 436160 516566 436172
rect 525794 436160 525800 436172
rect 525852 436160 525858 436212
rect 379146 436132 379152 436144
rect 378888 436104 379152 436132
rect 371694 436024 371700 436076
rect 371752 436064 371758 436076
rect 378888 436064 378916 436104
rect 379146 436092 379152 436104
rect 379204 436132 379210 436144
rect 395338 436132 395344 436144
rect 379204 436104 395344 436132
rect 379204 436092 379210 436104
rect 395338 436092 395344 436104
rect 395396 436092 395402 436144
rect 516134 436092 516140 436144
rect 516192 436132 516198 436144
rect 527174 436132 527180 436144
rect 516192 436104 527180 436132
rect 516192 436092 516198 436104
rect 527174 436092 527180 436104
rect 527232 436092 527238 436144
rect 371752 436036 378916 436064
rect 371752 436024 371758 436036
rect 371602 435956 371608 436008
rect 371660 435996 371666 436008
rect 378778 435996 378784 436008
rect 371660 435968 378784 435996
rect 371660 435956 371666 435968
rect 378778 435956 378784 435968
rect 378836 435996 378842 436008
rect 382918 435996 382924 436008
rect 378836 435968 382924 435996
rect 378836 435956 378842 435968
rect 382918 435956 382924 435968
rect 382976 435956 382982 436008
rect 516134 434800 516140 434852
rect 516192 434840 516198 434852
rect 521654 434840 521660 434852
rect 516192 434812 521660 434840
rect 516192 434800 516198 434812
rect 521654 434800 521660 434812
rect 521712 434800 521718 434852
rect 379054 434772 379060 434784
rect 378888 434744 379060 434772
rect 371694 434664 371700 434716
rect 371752 434704 371758 434716
rect 378888 434704 378916 434744
rect 379054 434732 379060 434744
rect 379112 434772 379118 434784
rect 393958 434772 393964 434784
rect 379112 434744 393964 434772
rect 379112 434732 379118 434744
rect 393958 434732 393964 434744
rect 394016 434732 394022 434784
rect 516226 434732 516232 434784
rect 516284 434772 516290 434784
rect 530026 434772 530032 434784
rect 516284 434744 530032 434772
rect 516284 434732 516290 434744
rect 530026 434732 530032 434744
rect 530084 434732 530090 434784
rect 371752 434676 378916 434704
rect 371752 434664 371758 434676
rect 371786 434596 371792 434648
rect 371844 434636 371850 434648
rect 376754 434636 376760 434648
rect 371844 434608 376760 434636
rect 371844 434596 371850 434608
rect 376754 434596 376760 434608
rect 376812 434636 376818 434648
rect 380158 434636 380164 434648
rect 376812 434608 380164 434636
rect 376812 434596 376818 434608
rect 380158 434596 380164 434608
rect 380216 434596 380222 434648
rect 371602 434528 371608 434580
rect 371660 434568 371666 434580
rect 375466 434568 375472 434580
rect 371660 434540 375472 434568
rect 371660 434528 371666 434540
rect 375466 434528 375472 434540
rect 375524 434568 375530 434580
rect 381538 434568 381544 434580
rect 375524 434540 381544 434568
rect 375524 434528 375530 434540
rect 381538 434528 381544 434540
rect 381596 434528 381602 434580
rect 444466 434392 444472 434444
rect 444524 434432 444530 434444
rect 446122 434432 446128 434444
rect 444524 434404 446128 434432
rect 444524 434392 444530 434404
rect 446122 434392 446128 434404
rect 446180 434392 446186 434444
rect 446122 433712 446128 433764
rect 446180 433752 446186 433764
rect 446858 433752 446864 433764
rect 446180 433724 446864 433752
rect 446180 433712 446186 433724
rect 446858 433712 446864 433724
rect 446916 433712 446922 433764
rect 516134 433440 516140 433492
rect 516192 433480 516198 433492
rect 524506 433480 524512 433492
rect 516192 433452 524512 433480
rect 516192 433440 516198 433452
rect 524506 433440 524512 433452
rect 524564 433440 524570 433492
rect 516502 433372 516508 433424
rect 516560 433412 516566 433424
rect 528646 433412 528652 433424
rect 516560 433384 528652 433412
rect 516560 433372 516566 433384
rect 528646 433372 528652 433384
rect 528704 433372 528710 433424
rect 516226 433304 516232 433356
rect 516284 433344 516290 433356
rect 530118 433344 530124 433356
rect 516284 433316 530124 433344
rect 516284 433304 516290 433316
rect 530118 433304 530124 433316
rect 530176 433304 530182 433356
rect 372154 433236 372160 433288
rect 372212 433276 372218 433288
rect 377490 433276 377496 433288
rect 372212 433248 377496 433276
rect 372212 433236 372218 433248
rect 377490 433236 377496 433248
rect 377548 433236 377554 433288
rect 444466 432896 444472 432948
rect 444524 432936 444530 432948
rect 446214 432936 446220 432948
rect 444524 432908 446220 432936
rect 444524 432896 444530 432908
rect 446214 432896 446220 432908
rect 446272 432936 446278 432948
rect 446766 432936 446772 432948
rect 446272 432908 446772 432936
rect 446272 432896 446278 432908
rect 446766 432896 446772 432908
rect 446824 432896 446830 432948
rect 376938 432800 376944 432812
rect 373966 432772 376944 432800
rect 371602 432624 371608 432676
rect 371660 432664 371666 432676
rect 373966 432664 373994 432772
rect 376938 432760 376944 432772
rect 376996 432800 377002 432812
rect 377398 432800 377404 432812
rect 376996 432772 377404 432800
rect 376996 432760 377002 432772
rect 377398 432760 377404 432772
rect 377456 432760 377462 432812
rect 371660 432636 373994 432664
rect 371660 432624 371666 432636
rect 378134 432624 378140 432676
rect 378192 432664 378198 432676
rect 378778 432664 378784 432676
rect 378192 432636 378784 432664
rect 378192 432624 378198 432636
rect 378778 432624 378784 432636
rect 378836 432624 378842 432676
rect 371694 432556 371700 432608
rect 371752 432596 371758 432608
rect 378152 432596 378180 432624
rect 371752 432568 378180 432596
rect 371752 432556 371758 432568
rect 371418 432420 371424 432472
rect 371476 432460 371482 432472
rect 371694 432460 371700 432472
rect 371476 432432 371700 432460
rect 371476 432420 371482 432432
rect 371694 432420 371700 432432
rect 371752 432420 371758 432472
rect 371326 432352 371332 432404
rect 371384 432352 371390 432404
rect 371344 432200 371372 432352
rect 371326 432148 371332 432200
rect 371384 432148 371390 432200
rect 371602 432148 371608 432200
rect 371660 432188 371666 432200
rect 372154 432188 372160 432200
rect 371660 432160 372160 432188
rect 371660 432148 371666 432160
rect 372154 432148 372160 432160
rect 372212 432148 372218 432200
rect 372154 432012 372160 432064
rect 372212 432052 372218 432064
rect 372430 432052 372436 432064
rect 372212 432024 372436 432052
rect 372212 432012 372218 432024
rect 372430 432012 372436 432024
rect 372488 432012 372494 432064
rect 516502 432012 516508 432064
rect 516560 432052 516566 432064
rect 525886 432052 525892 432064
rect 516560 432024 525892 432052
rect 516560 432012 516566 432024
rect 525886 432012 525892 432024
rect 525944 432012 525950 432064
rect 516778 431944 516784 431996
rect 516836 431984 516842 431996
rect 528554 431984 528560 431996
rect 516836 431956 528560 431984
rect 516836 431944 516842 431956
rect 528554 431944 528560 431956
rect 528612 431944 528618 431996
rect 443086 431060 443092 431112
rect 443144 431100 443150 431112
rect 446950 431100 446956 431112
rect 443144 431072 446956 431100
rect 443144 431060 443150 431072
rect 446950 431060 446956 431072
rect 447008 431060 447014 431112
rect 372062 429156 372068 429208
rect 372120 429196 372126 429208
rect 372522 429196 372528 429208
rect 372120 429168 372528 429196
rect 372120 429156 372126 429168
rect 372522 429156 372528 429168
rect 372580 429156 372586 429208
rect 371602 427048 371608 427100
rect 371660 427088 371666 427100
rect 376846 427088 376852 427100
rect 371660 427060 376852 427088
rect 371660 427048 371666 427060
rect 376846 427048 376852 427060
rect 376904 427048 376910 427100
rect 445570 426844 445576 426896
rect 445628 426884 445634 426896
rect 447410 426884 447416 426896
rect 445628 426856 447416 426884
rect 445628 426844 445634 426856
rect 447410 426844 447416 426856
rect 447468 426884 447474 426896
rect 447962 426884 447968 426896
rect 447468 426856 447968 426884
rect 447468 426844 447474 426856
rect 447962 426844 447968 426856
rect 448020 426844 448026 426896
rect 371602 426572 371608 426624
rect 371660 426612 371666 426624
rect 375834 426612 375840 426624
rect 371660 426584 375840 426612
rect 371660 426572 371666 426584
rect 375834 426572 375840 426584
rect 375892 426612 375898 426624
rect 376110 426612 376116 426624
rect 375892 426584 376116 426612
rect 375892 426572 375898 426584
rect 376110 426572 376116 426584
rect 376168 426572 376174 426624
rect 369118 426368 369124 426420
rect 369176 426408 369182 426420
rect 369486 426408 369492 426420
rect 369176 426380 369492 426408
rect 369176 426368 369182 426380
rect 369486 426368 369492 426380
rect 369544 426368 369550 426420
rect 371234 426368 371240 426420
rect 371292 426408 371298 426420
rect 375374 426408 375380 426420
rect 371292 426380 375380 426408
rect 371292 426368 371298 426380
rect 375374 426368 375380 426380
rect 375432 426368 375438 426420
rect 371602 426028 371608 426080
rect 371660 426068 371666 426080
rect 375466 426068 375472 426080
rect 371660 426040 375472 426068
rect 371660 426028 371666 426040
rect 375466 426028 375472 426040
rect 375524 426068 375530 426080
rect 376018 426068 376024 426080
rect 375524 426040 376024 426068
rect 375524 426028 375530 426040
rect 376018 426028 376024 426040
rect 376076 426028 376082 426080
rect 516778 425688 516784 425740
rect 516836 425728 516842 425740
rect 518158 425728 518164 425740
rect 516836 425700 518164 425728
rect 516836 425688 516842 425700
rect 518158 425688 518164 425700
rect 518216 425728 518222 425740
rect 524782 425728 524788 425740
rect 518216 425700 524788 425728
rect 518216 425688 518222 425700
rect 524782 425688 524788 425700
rect 524840 425688 524846 425740
rect 372614 425008 372620 425060
rect 372672 425048 372678 425060
rect 372982 425048 372988 425060
rect 372672 425020 372988 425048
rect 372672 425008 372678 425020
rect 372982 425008 372988 425020
rect 373040 425008 373046 425060
rect 371050 424668 371056 424720
rect 371108 424708 371114 424720
rect 374730 424708 374736 424720
rect 371108 424680 374736 424708
rect 371108 424668 371114 424680
rect 374730 424668 374736 424680
rect 374788 424668 374794 424720
rect 516134 424532 516140 424584
rect 516192 424572 516198 424584
rect 517790 424572 517796 424584
rect 516192 424544 517796 424572
rect 516192 424532 516198 424544
rect 517790 424532 517796 424544
rect 517848 424532 517854 424584
rect 516134 424396 516140 424448
rect 516192 424436 516198 424448
rect 518894 424436 518900 424448
rect 516192 424408 518900 424436
rect 516192 424396 516198 424408
rect 518894 424396 518900 424408
rect 518952 424436 518958 424448
rect 520458 424436 520464 424448
rect 518952 424408 520464 424436
rect 518952 424396 518958 424408
rect 520458 424396 520464 424408
rect 520516 424396 520522 424448
rect 516226 424328 516232 424380
rect 516284 424368 516290 424380
rect 522022 424368 522028 424380
rect 516284 424340 522028 424368
rect 516284 424328 516290 424340
rect 522022 424328 522028 424340
rect 522080 424328 522086 424380
rect 371602 423784 371608 423836
rect 371660 423824 371666 423836
rect 374914 423824 374920 423836
rect 371660 423796 374920 423824
rect 371660 423784 371666 423796
rect 374914 423784 374920 423796
rect 374972 423784 374978 423836
rect 371602 423648 371608 423700
rect 371660 423688 371666 423700
rect 371970 423688 371976 423700
rect 371660 423660 371976 423688
rect 371660 423648 371666 423660
rect 371970 423648 371976 423660
rect 372028 423648 372034 423700
rect 519170 423580 519176 423632
rect 519228 423620 519234 423632
rect 520642 423620 520648 423632
rect 519228 423592 520648 423620
rect 519228 423580 519234 423592
rect 520642 423580 520648 423592
rect 520700 423580 520706 423632
rect 371234 422560 371240 422612
rect 371292 422600 371298 422612
rect 374638 422600 374644 422612
rect 371292 422572 374644 422600
rect 371292 422560 371298 422572
rect 374638 422560 374644 422572
rect 374696 422560 374702 422612
rect 516134 422492 516140 422544
rect 516192 422532 516198 422544
rect 519170 422532 519176 422544
rect 516192 422504 519176 422532
rect 516192 422492 516198 422504
rect 519170 422492 519176 422504
rect 519228 422492 519234 422544
rect 516410 422464 516416 422476
rect 516152 422436 516416 422464
rect 516152 422408 516180 422436
rect 516410 422424 516416 422436
rect 516468 422424 516474 422476
rect 516134 422356 516140 422408
rect 516192 422356 516198 422408
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 273346 422328 273352 422340
rect 3476 422300 273352 422328
rect 3476 422288 3482 422300
rect 273346 422288 273352 422300
rect 273404 422288 273410 422340
rect 516318 422288 516324 422340
rect 516376 422328 516382 422340
rect 521930 422328 521936 422340
rect 516376 422300 521936 422328
rect 516376 422288 516382 422300
rect 521930 422288 521936 422300
rect 521988 422288 521994 422340
rect 516318 421880 516324 421932
rect 516376 421920 516382 421932
rect 517882 421920 517888 421932
rect 516376 421892 517888 421920
rect 516376 421880 516382 421892
rect 517882 421880 517888 421892
rect 517940 421880 517946 421932
rect 371142 421608 371148 421660
rect 371200 421648 371206 421660
rect 375006 421648 375012 421660
rect 371200 421620 375012 421648
rect 371200 421608 371206 421620
rect 375006 421608 375012 421620
rect 375064 421608 375070 421660
rect 371970 421540 371976 421592
rect 372028 421580 372034 421592
rect 374086 421580 374092 421592
rect 372028 421552 374092 421580
rect 372028 421540 372034 421552
rect 374086 421540 374092 421552
rect 374144 421580 374150 421592
rect 374822 421580 374828 421592
rect 374144 421552 374828 421580
rect 374144 421540 374150 421552
rect 374822 421540 374828 421552
rect 374880 421540 374886 421592
rect 516318 421540 516324 421592
rect 516376 421580 516382 421592
rect 520366 421580 520372 421592
rect 516376 421552 520372 421580
rect 516376 421540 516382 421552
rect 520366 421540 520372 421552
rect 520424 421540 520430 421592
rect 516318 421132 516324 421184
rect 516376 421172 516382 421184
rect 520642 421172 520648 421184
rect 516376 421144 520648 421172
rect 516376 421132 516382 421144
rect 520642 421132 520648 421144
rect 520700 421132 520706 421184
rect 446490 420928 446496 420980
rect 446548 420968 446554 420980
rect 449434 420968 449440 420980
rect 446548 420940 449440 420968
rect 446548 420928 446554 420940
rect 449434 420928 449440 420940
rect 449492 420928 449498 420980
rect 520366 420928 520372 420980
rect 520424 420968 520430 420980
rect 521746 420968 521752 420980
rect 520424 420940 521752 420968
rect 520424 420928 520430 420940
rect 521746 420928 521752 420940
rect 521804 420928 521810 420980
rect 443822 420860 443828 420912
rect 443880 420900 443886 420912
rect 449342 420900 449348 420912
rect 443880 420872 449348 420900
rect 443880 420860 443886 420872
rect 449342 420860 449348 420872
rect 449400 420860 449406 420912
rect 371970 420724 371976 420776
rect 372028 420764 372034 420776
rect 374270 420764 374276 420776
rect 372028 420736 374276 420764
rect 372028 420724 372034 420736
rect 374270 420724 374276 420736
rect 374328 420724 374334 420776
rect 445570 420588 445576 420640
rect 445628 420628 445634 420640
rect 446490 420628 446496 420640
rect 445628 420600 446496 420628
rect 445628 420588 445634 420600
rect 446490 420588 446496 420600
rect 446548 420588 446554 420640
rect 516778 420180 516784 420232
rect 516836 420220 516842 420232
rect 518250 420220 518256 420232
rect 516836 420192 518256 420220
rect 516836 420180 516842 420192
rect 518250 420180 518256 420192
rect 518308 420220 518314 420232
rect 520274 420220 520280 420232
rect 518308 420192 520280 420220
rect 518308 420180 518314 420192
rect 520274 420180 520280 420192
rect 520332 420180 520338 420232
rect 516778 419976 516784 420028
rect 516836 420016 516842 420028
rect 518066 420016 518072 420028
rect 516836 419988 518072 420016
rect 516836 419976 516842 419988
rect 518066 419976 518072 419988
rect 518124 420016 518130 420028
rect 518986 420016 518992 420028
rect 518124 419988 518992 420016
rect 518124 419976 518130 419988
rect 518986 419976 518992 419988
rect 519044 419976 519050 420028
rect 372430 419772 372436 419824
rect 372488 419812 372494 419824
rect 373902 419812 373908 419824
rect 372488 419784 373908 419812
rect 372488 419772 372494 419784
rect 373902 419772 373908 419784
rect 373960 419812 373966 419824
rect 374178 419812 374184 419824
rect 373960 419784 374184 419812
rect 373960 419772 373966 419784
rect 374178 419772 374184 419784
rect 374236 419772 374242 419824
rect 516318 419772 516324 419824
rect 516376 419812 516382 419824
rect 518894 419812 518900 419824
rect 516376 419784 518900 419812
rect 516376 419772 516382 419784
rect 518894 419772 518900 419784
rect 518952 419772 518958 419824
rect 373350 419432 373356 419484
rect 373408 419472 373414 419484
rect 374270 419472 374276 419484
rect 373408 419444 374276 419472
rect 373408 419432 373414 419444
rect 374270 419432 374276 419444
rect 374328 419432 374334 419484
rect 444466 419432 444472 419484
rect 444524 419472 444530 419484
rect 448698 419472 448704 419484
rect 444524 419444 448704 419472
rect 444524 419432 444530 419444
rect 448698 419432 448704 419444
rect 448756 419432 448762 419484
rect 371970 419092 371976 419144
rect 372028 419132 372034 419144
rect 374270 419132 374276 419144
rect 372028 419104 374276 419132
rect 372028 419092 372034 419104
rect 374270 419092 374276 419104
rect 374328 419092 374334 419144
rect 516502 418548 516508 418600
rect 516560 418588 516566 418600
rect 518986 418588 518992 418600
rect 516560 418560 518992 418588
rect 516560 418548 516566 418560
rect 518986 418548 518992 418560
rect 519044 418548 519050 418600
rect 516318 418480 516324 418532
rect 516376 418520 516382 418532
rect 519078 418520 519084 418532
rect 516376 418492 519084 418520
rect 516376 418480 516382 418492
rect 519078 418480 519084 418492
rect 519136 418480 519142 418532
rect 372154 418140 372160 418192
rect 372212 418180 372218 418192
rect 374454 418180 374460 418192
rect 372212 418152 374460 418180
rect 372212 418140 372218 418152
rect 373276 418124 373304 418152
rect 374454 418140 374460 418152
rect 374512 418140 374518 418192
rect 373258 418072 373264 418124
rect 373316 418072 373322 418124
rect 371970 417392 371976 417444
rect 372028 417432 372034 417444
rect 377306 417432 377312 417444
rect 372028 417404 377312 417432
rect 372028 417392 372034 417404
rect 377306 417392 377312 417404
rect 377364 417392 377370 417444
rect 516318 417392 516324 417444
rect 516376 417432 516382 417444
rect 517974 417432 517980 417444
rect 516376 417404 517980 417432
rect 516376 417392 516382 417404
rect 517974 417392 517980 417404
rect 518032 417392 518038 417444
rect 523126 417432 523132 417444
rect 518866 417404 523132 417432
rect 516594 417324 516600 417376
rect 516652 417364 516658 417376
rect 517698 417364 517704 417376
rect 516652 417336 517704 417364
rect 516652 417324 516658 417336
rect 517698 417324 517704 417336
rect 517756 417364 517762 417376
rect 518866 417364 518894 417404
rect 523126 417392 523132 417404
rect 523184 417392 523190 417444
rect 517756 417336 518894 417364
rect 517756 417324 517762 417336
rect 444650 417120 444656 417172
rect 444708 417160 444714 417172
rect 445846 417160 445852 417172
rect 444708 417132 445852 417160
rect 444708 417120 444714 417132
rect 445846 417120 445852 417132
rect 445904 417160 445910 417172
rect 446490 417160 446496 417172
rect 445904 417132 446496 417160
rect 445904 417120 445910 417132
rect 446490 417120 446496 417132
rect 446548 417120 446554 417172
rect 371970 416372 371976 416424
rect 372028 416412 372034 416424
rect 375558 416412 375564 416424
rect 372028 416384 375564 416412
rect 372028 416372 372034 416384
rect 375558 416372 375564 416384
rect 375616 416372 375622 416424
rect 516318 415760 516324 415812
rect 516376 415800 516382 415812
rect 520550 415800 520556 415812
rect 516376 415772 520556 415800
rect 516376 415760 516382 415772
rect 520550 415760 520556 415772
rect 520608 415760 520614 415812
rect 371970 415624 371976 415676
rect 372028 415664 372034 415676
rect 376018 415664 376024 415676
rect 372028 415636 376024 415664
rect 372028 415624 372034 415636
rect 376018 415624 376024 415636
rect 376076 415664 376082 415676
rect 377122 415664 377128 415676
rect 376076 415636 377128 415664
rect 376076 415624 376082 415636
rect 377122 415624 377128 415636
rect 377180 415624 377186 415676
rect 516502 415420 516508 415472
rect 516560 415460 516566 415472
rect 525978 415460 525984 415472
rect 516560 415432 525984 415460
rect 516560 415420 516566 415432
rect 525978 415420 525984 415432
rect 526036 415420 526042 415472
rect 444190 414808 444196 414860
rect 444248 414848 444254 414860
rect 447594 414848 447600 414860
rect 444248 414820 447600 414848
rect 444248 414808 444254 414820
rect 447594 414808 447600 414820
rect 447652 414808 447658 414860
rect 371970 414740 371976 414792
rect 372028 414780 372034 414792
rect 374546 414780 374552 414792
rect 372028 414752 374552 414780
rect 372028 414740 372034 414752
rect 374546 414740 374552 414752
rect 374604 414740 374610 414792
rect 516318 414672 516324 414724
rect 516376 414712 516382 414724
rect 519538 414712 519544 414724
rect 516376 414684 519544 414712
rect 516376 414672 516382 414684
rect 519538 414672 519544 414684
rect 519596 414712 519602 414724
rect 522114 414712 522120 414724
rect 519596 414684 522120 414712
rect 519596 414672 519602 414684
rect 522114 414672 522120 414684
rect 522172 414672 522178 414724
rect 516318 414060 516324 414112
rect 516376 414100 516382 414112
rect 523218 414100 523224 414112
rect 516376 414072 523224 414100
rect 516376 414060 516382 414072
rect 523218 414060 523224 414072
rect 523276 414060 523282 414112
rect 371234 413992 371240 414044
rect 371292 414032 371298 414044
rect 371292 414004 376156 414032
rect 371292 413992 371298 414004
rect 376128 413976 376156 414004
rect 516502 413992 516508 414044
rect 516560 414032 516566 414044
rect 524598 414032 524604 414044
rect 516560 414004 524604 414032
rect 516560 413992 516566 414004
rect 524598 413992 524604 414004
rect 524656 413992 524662 414044
rect 376110 413924 376116 413976
rect 376168 413964 376174 413976
rect 377214 413964 377220 413976
rect 376168 413936 377220 413964
rect 376168 413924 376174 413936
rect 377214 413924 377220 413936
rect 377272 413924 377278 413976
rect 445478 413652 445484 413704
rect 445536 413692 445542 413704
rect 447318 413692 447324 413704
rect 445536 413664 447324 413692
rect 445536 413652 445542 413664
rect 447318 413652 447324 413664
rect 447376 413652 447382 413704
rect 516318 413244 516324 413296
rect 516376 413284 516382 413296
rect 520918 413284 520924 413296
rect 516376 413256 520924 413284
rect 516376 413244 516382 413256
rect 520918 413244 520924 413256
rect 520976 413284 520982 413296
rect 524690 413284 524696 413296
rect 520976 413256 524696 413284
rect 520976 413244 520982 413256
rect 524690 413244 524696 413256
rect 524748 413244 524754 413296
rect 516778 412632 516784 412684
rect 516836 412672 516842 412684
rect 521838 412672 521844 412684
rect 516836 412644 521844 412672
rect 516836 412632 516842 412644
rect 521838 412632 521844 412644
rect 521896 412632 521902 412684
rect 445478 412564 445484 412616
rect 445536 412604 445542 412616
rect 447686 412604 447692 412616
rect 445536 412576 447692 412604
rect 445536 412564 445542 412576
rect 447686 412564 447692 412576
rect 447744 412564 447750 412616
rect 449250 412564 449256 412616
rect 449308 412604 449314 412616
rect 516226 412604 516232 412616
rect 449308 412576 516232 412604
rect 449308 412564 449314 412576
rect 516226 412564 516232 412576
rect 516284 412564 516290 412616
rect 372062 412496 372068 412548
rect 372120 412536 372126 412548
rect 372890 412536 372896 412548
rect 372120 412508 372896 412536
rect 372120 412496 372126 412508
rect 372890 412496 372896 412508
rect 372948 412496 372954 412548
rect 516318 412496 516324 412548
rect 516376 412536 516382 412548
rect 520366 412536 520372 412548
rect 516376 412508 520372 412536
rect 516376 412496 516382 412508
rect 520366 412496 520372 412508
rect 520424 412496 520430 412548
rect 371234 412088 371240 412140
rect 371292 412128 371298 412140
rect 375650 412128 375656 412140
rect 371292 412100 375656 412128
rect 371292 412088 371298 412100
rect 375650 412088 375656 412100
rect 375708 412088 375714 412140
rect 369118 412020 369124 412072
rect 369176 412060 369182 412072
rect 369762 412060 369768 412072
rect 369176 412032 369768 412060
rect 369176 412020 369182 412032
rect 369762 412020 369768 412032
rect 369820 412020 369826 412072
rect 500218 412020 500224 412072
rect 500276 412060 500282 412072
rect 516134 412060 516140 412072
rect 500276 412032 516140 412060
rect 500276 412020 500282 412032
rect 516134 412020 516140 412032
rect 516192 412020 516198 412072
rect 447686 411952 447692 412004
rect 447744 411992 447750 412004
rect 472710 411992 472716 412004
rect 447744 411964 472716 411992
rect 447744 411952 447750 411964
rect 472710 411952 472716 411964
rect 472768 411952 472774 412004
rect 497458 411952 497464 412004
rect 497516 411992 497522 412004
rect 516410 411992 516416 412004
rect 497516 411964 516416 411992
rect 497516 411952 497522 411964
rect 516410 411952 516416 411964
rect 516468 411952 516474 412004
rect 458818 411884 458824 411936
rect 458876 411924 458882 411936
rect 516502 411924 516508 411936
rect 458876 411896 516508 411924
rect 458876 411884 458882 411896
rect 516502 411884 516508 411896
rect 516560 411884 516566 411936
rect 472710 411272 472716 411324
rect 472768 411312 472774 411324
rect 513374 411312 513380 411324
rect 472768 411284 513380 411312
rect 472768 411272 472774 411284
rect 513374 411272 513380 411284
rect 513432 411272 513438 411324
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 274634 409884 274640 409896
rect 3200 409856 274640 409884
rect 3200 409844 3206 409856
rect 274634 409844 274640 409856
rect 274692 409844 274698 409896
rect 436830 409776 436836 409828
rect 436888 409816 436894 409828
rect 508958 409816 508964 409828
rect 436888 409788 508964 409816
rect 436888 409776 436894 409788
rect 508958 409776 508964 409788
rect 509016 409776 509022 409828
rect 432874 409708 432880 409760
rect 432932 409748 432938 409760
rect 504542 409748 504548 409760
rect 432932 409720 504548 409748
rect 432932 409708 432938 409720
rect 504542 409708 504548 409720
rect 504600 409708 504606 409760
rect 441062 409640 441068 409692
rect 441120 409680 441126 409692
rect 513006 409680 513012 409692
rect 441120 409652 513012 409680
rect 441120 409640 441126 409652
rect 513006 409640 513012 409652
rect 513064 409640 513070 409692
rect 304258 409164 304264 409216
rect 304316 409204 304322 409216
rect 366910 409204 366916 409216
rect 304316 409176 366916 409204
rect 304316 409164 304322 409176
rect 366910 409164 366916 409176
rect 366968 409164 366974 409216
rect 304350 409096 304356 409148
rect 304408 409136 304414 409148
rect 438854 409136 438860 409148
rect 304408 409108 438860 409136
rect 304408 409096 304414 409108
rect 438854 409096 438860 409108
rect 438912 409096 438918 409148
rect 501598 409096 501604 409148
rect 501656 409136 501662 409148
rect 510982 409136 510988 409148
rect 501656 409108 510988 409136
rect 501656 409096 501662 409108
rect 510982 409096 510988 409108
rect 511040 409096 511046 409148
rect 431954 408484 431960 408536
rect 432012 408524 432018 408536
rect 432874 408524 432880 408536
rect 432012 408496 432880 408524
rect 432012 408484 432018 408496
rect 432874 408484 432880 408496
rect 432932 408484 432938 408536
rect 223390 404336 223396 404388
rect 223448 404376 223454 404388
rect 580166 404376 580172 404388
rect 223448 404348 580172 404376
rect 223448 404336 223454 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 387058 398080 387064 398132
rect 387116 398120 387122 398132
rect 450078 398120 450084 398132
rect 387116 398092 450084 398120
rect 387116 398080 387122 398092
rect 450078 398080 450084 398092
rect 450136 398080 450142 398132
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 274726 397508 274732 397520
rect 3476 397480 274732 397508
rect 3476 397468 3482 397480
rect 274726 397468 274732 397480
rect 274784 397468 274790 397520
rect 395338 395972 395344 396024
rect 395396 396012 395402 396024
rect 395982 396012 395988 396024
rect 395396 395984 395988 396012
rect 395396 395972 395402 395984
rect 395982 395972 395988 395984
rect 396040 395972 396046 396024
rect 395982 395292 395988 395344
rect 396040 395332 396046 395344
rect 449986 395332 449992 395344
rect 396040 395304 449992 395332
rect 396040 395292 396046 395304
rect 449986 395292 449992 395304
rect 450044 395292 450050 395344
rect 393958 394612 393964 394664
rect 394016 394652 394022 394664
rect 394602 394652 394608 394664
rect 394016 394624 394608 394652
rect 394016 394612 394022 394624
rect 394602 394612 394608 394624
rect 394660 394612 394666 394664
rect 394602 393932 394608 393984
rect 394660 393972 394666 393984
rect 450538 393972 450544 393984
rect 394660 393944 450544 393972
rect 394660 393932 394666 393944
rect 450538 393932 450544 393944
rect 450596 393932 450602 393984
rect 446858 389172 446864 389224
rect 446916 389212 446922 389224
rect 447410 389212 447416 389224
rect 446916 389184 447416 389212
rect 446916 389172 446922 389184
rect 447410 389172 447416 389184
rect 447468 389212 447474 389224
rect 517882 389212 517888 389224
rect 447468 389184 517888 389212
rect 447468 389172 447474 389184
rect 517882 389172 517888 389184
rect 517940 389172 517946 389224
rect 399478 388424 399484 388476
rect 399536 388464 399542 388476
rect 400122 388464 400128 388476
rect 399536 388436 400128 388464
rect 399536 388424 399542 388436
rect 400122 388424 400128 388436
rect 400180 388464 400186 388476
rect 448698 388464 448704 388476
rect 400180 388436 448704 388464
rect 400180 388424 400186 388436
rect 448698 388424 448704 388436
rect 448756 388464 448762 388476
rect 449158 388464 449164 388476
rect 448756 388436 449164 388464
rect 448756 388424 448762 388436
rect 449158 388424 449164 388436
rect 449216 388424 449222 388476
rect 382918 387064 382924 387116
rect 382976 387104 382982 387116
rect 383562 387104 383568 387116
rect 382976 387076 383568 387104
rect 382976 387064 382982 387076
rect 383562 387064 383568 387076
rect 383620 387104 383626 387116
rect 441706 387104 441712 387116
rect 383620 387076 441712 387104
rect 383620 387064 383626 387076
rect 441706 387064 441712 387076
rect 441764 387064 441770 387116
rect 377398 385636 377404 385688
rect 377456 385676 377462 385688
rect 448606 385676 448612 385688
rect 377456 385648 448612 385676
rect 377456 385636 377462 385648
rect 448606 385636 448612 385648
rect 448664 385636 448670 385688
rect 380158 384276 380164 384328
rect 380216 384316 380222 384328
rect 448514 384316 448520 384328
rect 380216 384288 448520 384316
rect 380216 384276 380222 384288
rect 448514 384276 448520 384288
rect 448572 384276 448578 384328
rect 446766 381488 446772 381540
rect 446824 381528 446830 381540
rect 520642 381528 520648 381540
rect 446824 381500 520648 381528
rect 446824 381488 446830 381500
rect 520642 381488 520648 381500
rect 520700 381488 520706 381540
rect 446490 380128 446496 380180
rect 446548 380168 446554 380180
rect 523218 380168 523224 380180
rect 446548 380140 523224 380168
rect 446548 380128 446554 380140
rect 523218 380128 523224 380140
rect 523276 380128 523282 380180
rect 446490 379516 446496 379568
rect 446548 379556 446554 379568
rect 447042 379556 447048 379568
rect 446548 379528 447048 379556
rect 446548 379516 446554 379528
rect 447042 379516 447048 379528
rect 447100 379516 447106 379568
rect 222102 378156 222108 378208
rect 222160 378196 222166 378208
rect 580166 378196 580172 378208
rect 222160 378168 580172 378196
rect 222160 378156 222166 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 446674 378088 446680 378140
rect 446732 378128 446738 378140
rect 447502 378128 447508 378140
rect 446732 378100 447508 378128
rect 446732 378088 446738 378100
rect 447502 378088 447508 378100
rect 447560 378088 447566 378140
rect 516594 377408 516600 377460
rect 516652 377448 516658 377460
rect 522022 377448 522028 377460
rect 516652 377420 522028 377448
rect 516652 377408 516658 377420
rect 522022 377408 522028 377420
rect 522080 377408 522086 377460
rect 447502 376728 447508 376780
rect 447560 376768 447566 376780
rect 516410 376768 516416 376780
rect 447560 376740 516416 376768
rect 447560 376728 447566 376740
rect 516410 376728 516416 376740
rect 516468 376768 516474 376780
rect 516594 376768 516600 376780
rect 516468 376740 516600 376768
rect 516468 376728 516474 376740
rect 516594 376728 516600 376740
rect 516652 376728 516658 376780
rect 447962 375980 447968 376032
rect 448020 376020 448026 376032
rect 519078 376020 519084 376032
rect 448020 375992 519084 376020
rect 448020 375980 448026 375992
rect 519078 375980 519084 375992
rect 519136 375980 519142 376032
rect 449342 373260 449348 373312
rect 449400 373300 449406 373312
rect 520550 373300 520556 373312
rect 449400 373272 520556 373300
rect 449400 373260 449406 373272
rect 520550 373260 520556 373272
rect 520608 373260 520614 373312
rect 378778 371832 378784 371884
rect 378836 371872 378842 371884
rect 441614 371872 441620 371884
rect 378836 371844 441620 371872
rect 378836 371832 378842 371844
rect 441614 371832 441620 371844
rect 441672 371832 441678 371884
rect 516134 371696 516140 371748
rect 516192 371736 516198 371748
rect 519170 371736 519176 371748
rect 516192 371708 519176 371736
rect 516192 371696 516198 371708
rect 519170 371696 519176 371708
rect 519228 371696 519234 371748
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 276014 371260 276020 371272
rect 3476 371232 276020 371260
rect 3476 371220 3482 371232
rect 276014 371220 276020 371232
rect 276072 371220 276078 371272
rect 446490 371220 446496 371272
rect 446548 371260 446554 371272
rect 516134 371260 516140 371272
rect 446548 371232 516140 371260
rect 446548 371220 446554 371232
rect 516134 371220 516140 371232
rect 516192 371220 516198 371272
rect 506474 370472 506480 370524
rect 506532 370512 506538 370524
rect 513374 370512 513380 370524
rect 506532 370484 513380 370512
rect 506532 370472 506538 370484
rect 513374 370472 513380 370484
rect 513432 370472 513438 370524
rect 381538 369860 381544 369912
rect 381596 369900 381602 369912
rect 382182 369900 382188 369912
rect 381596 369872 382188 369900
rect 381596 369860 381602 369872
rect 382182 369860 382188 369872
rect 382240 369900 382246 369912
rect 444466 369900 444472 369912
rect 382240 369872 444472 369900
rect 382240 369860 382246 369872
rect 444466 369860 444472 369872
rect 444524 369900 444530 369912
rect 449894 369900 449900 369912
rect 444524 369872 449900 369900
rect 444524 369860 444530 369872
rect 449894 369860 449900 369872
rect 449952 369860 449958 369912
rect 516134 369792 516140 369844
rect 516192 369832 516198 369844
rect 524782 369832 524788 369844
rect 516192 369804 524788 369832
rect 516192 369792 516198 369804
rect 524782 369792 524788 369804
rect 524840 369792 524846 369844
rect 372614 369656 372620 369708
rect 372672 369696 372678 369708
rect 372890 369696 372896 369708
rect 372672 369668 372896 369696
rect 372672 369656 372678 369668
rect 372890 369656 372896 369668
rect 372948 369656 372954 369708
rect 371786 369520 371792 369572
rect 371844 369560 371850 369572
rect 372614 369560 372620 369572
rect 371844 369532 372620 369560
rect 371844 369520 371850 369532
rect 372614 369520 372620 369532
rect 372672 369520 372678 369572
rect 370958 369316 370964 369368
rect 371016 369356 371022 369368
rect 374730 369356 374736 369368
rect 371016 369328 374736 369356
rect 371016 369316 371022 369328
rect 374730 369316 374736 369328
rect 374788 369356 374794 369368
rect 377582 369356 377588 369368
rect 374788 369328 377588 369356
rect 374788 369316 374794 369328
rect 377582 369316 377588 369328
rect 377640 369316 377646 369368
rect 373994 369248 374000 369300
rect 374052 369288 374058 369300
rect 441614 369288 441620 369300
rect 374052 369260 441620 369288
rect 374052 369248 374058 369260
rect 441614 369248 441620 369260
rect 441672 369248 441678 369300
rect 375282 369180 375288 369232
rect 375340 369220 375346 369232
rect 441338 369220 441344 369232
rect 375340 369192 441344 369220
rect 375340 369180 375346 369192
rect 441338 369180 441344 369192
rect 441396 369180 441402 369232
rect 372614 369112 372620 369164
rect 372672 369152 372678 369164
rect 442258 369152 442264 369164
rect 372672 369124 442264 369152
rect 372672 369112 372678 369124
rect 442258 369112 442264 369124
rect 442316 369112 442322 369164
rect 447870 369112 447876 369164
rect 447928 369152 447934 369164
rect 513742 369152 513748 369164
rect 447928 369124 513748 369152
rect 447928 369112 447934 369124
rect 513742 369112 513748 369124
rect 513800 369112 513806 369164
rect 371418 368500 371424 368552
rect 371476 368540 371482 368552
rect 375282 368540 375288 368552
rect 371476 368512 375288 368540
rect 371476 368500 371482 368512
rect 375282 368500 375288 368512
rect 375340 368500 375346 368552
rect 516134 368364 516140 368416
rect 516192 368404 516198 368416
rect 517790 368404 517796 368416
rect 516192 368376 517796 368404
rect 516192 368364 516198 368376
rect 517790 368364 517796 368376
rect 517848 368364 517854 368416
rect 389082 367888 389088 367940
rect 389140 367928 389146 367940
rect 441614 367928 441620 367940
rect 389140 367900 441620 367928
rect 389140 367888 389146 367900
rect 441614 367888 441620 367900
rect 441672 367888 441678 367940
rect 455322 367888 455328 367940
rect 455380 367928 455386 367940
rect 513650 367928 513656 367940
rect 455380 367900 513656 367928
rect 455380 367888 455386 367900
rect 513650 367888 513656 367900
rect 513708 367888 513714 367940
rect 390462 367820 390468 367872
rect 390520 367860 390526 367872
rect 441338 367860 441344 367872
rect 390520 367832 441344 367860
rect 390520 367820 390526 367832
rect 441338 367820 441344 367832
rect 441396 367860 441402 367872
rect 444558 367860 444564 367872
rect 441396 367832 444564 367860
rect 441396 367820 441402 367832
rect 444558 367820 444564 367832
rect 444616 367820 444622 367872
rect 502978 367820 502984 367872
rect 503036 367860 503042 367872
rect 513742 367860 513748 367872
rect 503036 367832 513748 367860
rect 503036 367820 503042 367832
rect 513742 367820 513748 367832
rect 513800 367820 513806 367872
rect 370590 367752 370596 367804
rect 370648 367792 370654 367804
rect 374638 367792 374644 367804
rect 370648 367764 374644 367792
rect 370648 367752 370654 367764
rect 374638 367752 374644 367764
rect 374696 367792 374702 367804
rect 377490 367792 377496 367804
rect 374696 367764 377496 367792
rect 374696 367752 374702 367764
rect 377490 367752 377496 367764
rect 377548 367752 377554 367804
rect 516134 367752 516140 367804
rect 516192 367792 516198 367804
rect 520458 367792 520464 367804
rect 516192 367764 520464 367792
rect 516192 367752 516198 367764
rect 520458 367752 520464 367764
rect 520516 367752 520522 367804
rect 370314 367480 370320 367532
rect 370372 367520 370378 367532
rect 372890 367520 372896 367532
rect 370372 367492 372896 367520
rect 370372 367480 370378 367492
rect 372890 367480 372896 367492
rect 372948 367480 372954 367532
rect 371326 367140 371332 367192
rect 371384 367180 371390 367192
rect 373994 367180 374000 367192
rect 371384 367152 374000 367180
rect 371384 367140 371390 367152
rect 373994 367140 374000 367152
rect 374052 367140 374058 367192
rect 444282 367004 444288 367056
rect 444340 367044 444346 367056
rect 444742 367044 444748 367056
rect 444340 367016 444748 367044
rect 444340 367004 444346 367016
rect 444742 367004 444748 367016
rect 444800 367004 444806 367056
rect 447778 366936 447784 366988
rect 447836 366976 447842 366988
rect 454034 366976 454040 366988
rect 447836 366948 454040 366976
rect 447836 366936 447842 366948
rect 454034 366936 454040 366948
rect 454092 366976 454098 366988
rect 455322 366976 455328 366988
rect 454092 366948 455328 366976
rect 454092 366936 454098 366948
rect 455322 366936 455328 366948
rect 455380 366936 455386 366988
rect 370958 366460 370964 366512
rect 371016 366500 371022 366512
rect 374914 366500 374920 366512
rect 371016 366472 374920 366500
rect 371016 366460 371022 366472
rect 374914 366460 374920 366472
rect 374972 366500 374978 366512
rect 377030 366500 377036 366512
rect 374972 366472 377036 366500
rect 374972 366460 374978 366472
rect 377030 366460 377036 366472
rect 377088 366460 377094 366512
rect 444650 365712 444656 365764
rect 444708 365752 444714 365764
rect 452654 365752 452660 365764
rect 444708 365724 452660 365752
rect 444708 365712 444714 365724
rect 452654 365712 452660 365724
rect 452712 365712 452718 365764
rect 444926 365644 444932 365696
rect 444984 365684 444990 365696
rect 448698 365684 448704 365696
rect 444984 365656 448704 365684
rect 444984 365644 444990 365656
rect 448698 365644 448704 365656
rect 448756 365644 448762 365696
rect 370958 364760 370964 364812
rect 371016 364800 371022 364812
rect 373994 364800 374000 364812
rect 371016 364772 374000 364800
rect 371016 364760 371022 364772
rect 373994 364760 374000 364772
rect 374052 364800 374058 364812
rect 375006 364800 375012 364812
rect 374052 364772 375012 364800
rect 374052 364760 374058 364772
rect 375006 364760 375012 364772
rect 375064 364760 375070 364812
rect 444190 364352 444196 364404
rect 444248 364392 444254 364404
rect 451274 364392 451280 364404
rect 444248 364364 451280 364392
rect 444248 364352 444254 364364
rect 451274 364352 451280 364364
rect 451332 364352 451338 364404
rect 445570 364284 445576 364336
rect 445628 364324 445634 364336
rect 450078 364324 450084 364336
rect 445628 364296 450084 364324
rect 445628 364284 445634 364296
rect 450078 364284 450084 364296
rect 450136 364284 450142 364336
rect 445110 363808 445116 363860
rect 445168 363848 445174 363860
rect 449986 363848 449992 363860
rect 445168 363820 449992 363848
rect 445168 363808 445174 363820
rect 449986 363808 449992 363820
rect 450044 363808 450050 363860
rect 516134 363604 516140 363656
rect 516192 363644 516198 363656
rect 521930 363644 521936 363656
rect 516192 363616 521936 363644
rect 516192 363604 516198 363616
rect 521930 363604 521936 363616
rect 521988 363604 521994 363656
rect 369118 363536 369124 363588
rect 369176 363576 369182 363588
rect 370314 363576 370320 363588
rect 369176 363548 370320 363576
rect 369176 363536 369182 363548
rect 370314 363536 370320 363548
rect 370372 363536 370378 363588
rect 386322 362924 386328 362976
rect 386380 362964 386386 362976
rect 387058 362964 387064 362976
rect 386380 362936 387064 362964
rect 386380 362924 386386 362936
rect 387058 362924 387064 362936
rect 387116 362924 387122 362976
rect 445110 362856 445116 362908
rect 445168 362896 445174 362908
rect 450170 362896 450176 362908
rect 445168 362868 450176 362896
rect 445168 362856 445174 362868
rect 450170 362856 450176 362868
rect 450228 362856 450234 362908
rect 516134 362652 516140 362704
rect 516192 362692 516198 362704
rect 517882 362692 517888 362704
rect 516192 362664 517888 362692
rect 516192 362652 516198 362664
rect 517882 362652 517888 362664
rect 517940 362652 517946 362704
rect 370958 362448 370964 362500
rect 371016 362488 371022 362500
rect 374086 362488 374092 362500
rect 371016 362460 374092 362488
rect 371016 362448 371022 362460
rect 374086 362448 374092 362460
rect 374144 362448 374150 362500
rect 445110 361496 445116 361548
rect 445168 361536 445174 361548
rect 448514 361536 448520 361548
rect 445168 361508 448520 361536
rect 445168 361496 445174 361508
rect 448514 361496 448520 361508
rect 448572 361496 448578 361548
rect 516778 360816 516784 360868
rect 516836 360856 516842 360868
rect 518250 360856 518256 360868
rect 516836 360828 518256 360856
rect 516836 360816 516842 360828
rect 518250 360816 518256 360828
rect 518308 360856 518314 360868
rect 521746 360856 521752 360868
rect 518308 360828 521752 360856
rect 518308 360816 518314 360828
rect 521746 360816 521752 360828
rect 521804 360816 521810 360868
rect 516134 360680 516140 360732
rect 516192 360720 516198 360732
rect 520642 360720 520648 360732
rect 516192 360692 520648 360720
rect 516192 360680 516198 360692
rect 520642 360680 520648 360692
rect 520700 360680 520706 360732
rect 378042 360204 378048 360256
rect 378100 360244 378106 360256
rect 378778 360244 378784 360256
rect 378100 360216 378784 360244
rect 378100 360204 378106 360216
rect 378778 360204 378784 360216
rect 378836 360204 378842 360256
rect 379422 360204 379428 360256
rect 379480 360244 379486 360256
rect 380158 360244 380164 360256
rect 379480 360216 380164 360244
rect 379480 360204 379486 360216
rect 380158 360204 380164 360216
rect 380216 360204 380222 360256
rect 445110 360136 445116 360188
rect 445168 360176 445174 360188
rect 448606 360176 448612 360188
rect 445168 360148 448612 360176
rect 445168 360136 445174 360148
rect 448606 360136 448612 360148
rect 448664 360136 448670 360188
rect 376662 359252 376668 359304
rect 376720 359292 376726 359304
rect 377398 359292 377404 359304
rect 376720 359264 377404 359292
rect 376720 359252 376726 359264
rect 377398 359252 377404 359264
rect 377456 359252 377462 359304
rect 369762 359116 369768 359168
rect 369820 359156 369826 359168
rect 373350 359156 373356 359168
rect 369820 359128 373356 359156
rect 369820 359116 369826 359128
rect 373350 359116 373356 359128
rect 373408 359116 373414 359168
rect 516134 359116 516140 359168
rect 516192 359156 516198 359168
rect 518894 359156 518900 359168
rect 516192 359128 518900 359156
rect 516192 359116 516198 359128
rect 518894 359116 518900 359128
rect 518952 359156 518958 359168
rect 519170 359156 519176 359168
rect 518952 359128 519176 359156
rect 518952 359116 518958 359128
rect 519170 359116 519176 359128
rect 519228 359116 519234 359168
rect 445662 358708 445668 358760
rect 445720 358748 445726 358760
rect 497458 358748 497464 358760
rect 445720 358720 497464 358748
rect 445720 358708 445726 358720
rect 497458 358708 497464 358720
rect 497516 358708 497522 358760
rect 516134 357892 516140 357944
rect 516192 357932 516198 357944
rect 520274 357932 520280 357944
rect 516192 357904 520280 357932
rect 516192 357892 516198 357904
rect 520274 357892 520280 357904
rect 520332 357892 520338 357944
rect 370682 357824 370688 357876
rect 370740 357864 370746 357876
rect 373350 357864 373356 357876
rect 370740 357836 373356 357864
rect 370740 357824 370746 357836
rect 373350 357824 373356 357836
rect 373408 357824 373414 357876
rect 369762 357756 369768 357808
rect 369820 357796 369826 357808
rect 370130 357796 370136 357808
rect 369820 357768 370136 357796
rect 369820 357756 369826 357768
rect 370130 357756 370136 357768
rect 370188 357756 370194 357808
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 277394 357456 277400 357468
rect 3200 357428 277400 357456
rect 3200 357416 3206 357428
rect 277394 357416 277400 357428
rect 277452 357416 277458 357468
rect 445570 357348 445576 357400
rect 445628 357388 445634 357400
rect 500218 357388 500224 357400
rect 445628 357360 500224 357388
rect 445628 357348 445634 357360
rect 500218 357348 500224 357360
rect 500276 357348 500282 357400
rect 516410 357348 516416 357400
rect 516468 357388 516474 357400
rect 518066 357388 518072 357400
rect 516468 357360 518072 357388
rect 516468 357348 516474 357360
rect 518066 357348 518072 357360
rect 518124 357348 518130 357400
rect 445478 357280 445484 357332
rect 445536 357320 445542 357332
rect 458818 357320 458824 357332
rect 445536 357292 458824 357320
rect 445536 357280 445542 357292
rect 458818 357280 458824 357292
rect 458876 357280 458882 357332
rect 370958 356736 370964 356788
rect 371016 356776 371022 356788
rect 374178 356776 374184 356788
rect 371016 356748 374184 356776
rect 371016 356736 371022 356748
rect 374178 356736 374184 356748
rect 374236 356736 374242 356788
rect 516134 355580 516140 355632
rect 516192 355620 516198 355632
rect 518986 355620 518992 355632
rect 516192 355592 518992 355620
rect 516192 355580 516198 355592
rect 518986 355580 518992 355592
rect 519044 355580 519050 355632
rect 370958 355512 370964 355564
rect 371016 355552 371022 355564
rect 374270 355552 374276 355564
rect 371016 355524 374276 355552
rect 371016 355512 371022 355524
rect 374270 355512 374276 355524
rect 374328 355512 374334 355564
rect 445018 355308 445024 355360
rect 445076 355348 445082 355360
rect 457438 355348 457444 355360
rect 445076 355320 457444 355348
rect 445076 355308 445082 355320
rect 457438 355308 457444 355320
rect 457496 355308 457502 355360
rect 516134 354492 516140 354544
rect 516192 354532 516198 354544
rect 519078 354532 519084 354544
rect 516192 354504 519084 354532
rect 516192 354492 516198 354504
rect 519078 354492 519084 354504
rect 519136 354492 519142 354544
rect 370958 354424 370964 354476
rect 371016 354464 371022 354476
rect 373258 354464 373264 354476
rect 371016 354436 373264 354464
rect 371016 354424 371022 354436
rect 373258 354424 373264 354436
rect 373316 354424 373322 354476
rect 445570 354016 445576 354068
rect 445628 354056 445634 354068
rect 448422 354056 448428 354068
rect 445628 354028 448428 354056
rect 445628 354016 445634 354028
rect 448422 354016 448428 354028
rect 448480 354056 448486 354068
rect 449250 354056 449256 354068
rect 448480 354028 449256 354056
rect 448480 354016 448486 354028
rect 449250 354016 449256 354028
rect 449308 354016 449314 354068
rect 445110 353812 445116 353864
rect 445168 353852 445174 353864
rect 446122 353852 446128 353864
rect 445168 353824 446128 353852
rect 445168 353812 445174 353824
rect 446122 353812 446128 353824
rect 446180 353852 446186 353864
rect 447870 353852 447876 353864
rect 446180 353824 447876 353852
rect 446180 353812 446186 353824
rect 447870 353812 447876 353824
rect 447928 353812 447934 353864
rect 446214 353336 446220 353388
rect 446272 353376 446278 353388
rect 447962 353376 447968 353388
rect 446272 353348 447968 353376
rect 446272 353336 446278 353348
rect 447962 353336 447968 353348
rect 448020 353336 448026 353388
rect 444650 353268 444656 353320
rect 444708 353308 444714 353320
rect 449158 353308 449164 353320
rect 444708 353280 449164 353308
rect 444708 353268 444714 353280
rect 449158 353268 449164 353280
rect 449216 353268 449222 353320
rect 445570 352588 445576 352640
rect 445628 352628 445634 352640
rect 446030 352628 446036 352640
rect 445628 352600 446036 352628
rect 445628 352588 445634 352600
rect 446030 352588 446036 352600
rect 446088 352628 446094 352640
rect 454034 352628 454040 352640
rect 446088 352600 454040 352628
rect 446088 352588 446094 352600
rect 454034 352588 454040 352600
rect 454092 352588 454098 352640
rect 502978 352560 502984 352572
rect 451246 352532 502984 352560
rect 445570 352452 445576 352504
rect 445628 352492 445634 352504
rect 447134 352492 447140 352504
rect 445628 352464 447140 352492
rect 445628 352452 445634 352464
rect 447134 352452 447140 352464
rect 447192 352492 447198 352504
rect 448606 352492 448612 352504
rect 447192 352464 448612 352492
rect 447192 352452 447198 352464
rect 448606 352452 448612 352464
rect 448664 352492 448670 352504
rect 451246 352492 451274 352532
rect 502978 352520 502984 352532
rect 503036 352520 503042 352572
rect 448664 352464 451274 352492
rect 448664 352452 448670 352464
rect 370866 352112 370872 352164
rect 370924 352152 370930 352164
rect 374362 352152 374368 352164
rect 370924 352124 374368 352152
rect 370924 352112 370930 352124
rect 374362 352112 374368 352124
rect 374420 352112 374426 352164
rect 445570 351908 445576 351960
rect 445628 351948 445634 351960
rect 447502 351948 447508 351960
rect 445628 351920 447508 351948
rect 445628 351908 445634 351920
rect 447502 351908 447508 351920
rect 447560 351908 447566 351960
rect 516134 351840 516140 351892
rect 516192 351880 516198 351892
rect 523126 351880 523132 351892
rect 516192 351852 523132 351880
rect 516192 351840 516198 351852
rect 523126 351840 523132 351852
rect 523184 351840 523190 351892
rect 444374 351364 444380 351416
rect 444432 351404 444438 351416
rect 446490 351404 446496 351416
rect 444432 351376 446496 351404
rect 444432 351364 444438 351376
rect 446490 351364 446496 351376
rect 446548 351364 446554 351416
rect 370682 351160 370688 351212
rect 370740 351200 370746 351212
rect 377122 351200 377128 351212
rect 370740 351172 377128 351200
rect 370740 351160 370746 351172
rect 377122 351160 377128 351172
rect 377180 351160 377186 351212
rect 370590 350888 370596 350940
rect 370648 350928 370654 350940
rect 372614 350928 372620 350940
rect 370648 350900 372620 350928
rect 370648 350888 370654 350900
rect 372614 350888 372620 350900
rect 372672 350888 372678 350940
rect 523126 350548 523132 350600
rect 523184 350588 523190 350600
rect 524782 350588 524788 350600
rect 523184 350560 524788 350588
rect 523184 350548 523190 350560
rect 524782 350548 524788 350560
rect 524840 350548 524846 350600
rect 443822 350480 443828 350532
rect 443880 350520 443886 350532
rect 444374 350520 444380 350532
rect 443880 350492 444380 350520
rect 443880 350480 443886 350492
rect 444374 350480 444380 350492
rect 444432 350480 444438 350532
rect 445478 350208 445484 350260
rect 445536 350248 445542 350260
rect 447410 350248 447416 350260
rect 445536 350220 447416 350248
rect 445536 350208 445542 350220
rect 447410 350208 447416 350220
rect 447468 350208 447474 350260
rect 370958 349800 370964 349852
rect 371016 349840 371022 349852
rect 375558 349840 375564 349852
rect 371016 349812 375564 349840
rect 371016 349800 371022 349812
rect 375558 349800 375564 349812
rect 375616 349840 375622 349852
rect 377214 349840 377220 349852
rect 375616 349812 377220 349840
rect 375616 349800 375622 349812
rect 377214 349800 377220 349812
rect 377272 349800 377278 349852
rect 516594 349800 516600 349852
rect 516652 349840 516658 349852
rect 517698 349840 517704 349852
rect 516652 349812 517704 349840
rect 516652 349800 516658 349812
rect 517698 349800 517704 349812
rect 517756 349840 517762 349852
rect 525978 349840 525984 349852
rect 517756 349812 525984 349840
rect 517756 349800 517762 349812
rect 525978 349800 525984 349812
rect 526036 349800 526042 349852
rect 445938 349664 445944 349716
rect 445996 349704 446002 349716
rect 446766 349704 446772 349716
rect 445996 349676 446772 349704
rect 445996 349664 446002 349676
rect 446766 349664 446772 349676
rect 446824 349664 446830 349716
rect 516134 348780 516140 348832
rect 516192 348820 516198 348832
rect 520550 348820 520556 348832
rect 516192 348792 520556 348820
rect 516192 348780 516198 348792
rect 520550 348780 520556 348792
rect 520608 348780 520614 348832
rect 370958 348644 370964 348696
rect 371016 348684 371022 348696
rect 376018 348684 376024 348696
rect 371016 348656 376024 348684
rect 371016 348644 371022 348656
rect 376018 348644 376024 348656
rect 376076 348644 376082 348696
rect 441890 347692 441896 347744
rect 441948 347732 441954 347744
rect 443270 347732 443276 347744
rect 441948 347704 443276 347732
rect 441948 347692 441954 347704
rect 443270 347692 443276 347704
rect 443328 347692 443334 347744
rect 445846 347692 445852 347744
rect 445904 347732 445910 347744
rect 446306 347732 446312 347744
rect 445904 347704 446312 347732
rect 445904 347692 445910 347704
rect 446306 347692 446312 347704
rect 446364 347692 446370 347744
rect 521010 347692 521016 347744
rect 521068 347732 521074 347744
rect 524598 347732 524604 347744
rect 521068 347704 524604 347732
rect 521068 347692 521074 347704
rect 524598 347692 524604 347704
rect 524656 347692 524662 347744
rect 370498 347148 370504 347200
rect 370556 347188 370562 347200
rect 375558 347188 375564 347200
rect 370556 347160 375564 347188
rect 370556 347148 370562 347160
rect 375558 347148 375564 347160
rect 375616 347188 375622 347200
rect 376110 347188 376116 347200
rect 375616 347160 376116 347188
rect 375616 347148 375622 347160
rect 376110 347148 376116 347160
rect 376168 347148 376174 347200
rect 516134 347012 516140 347064
rect 516192 347052 516198 347064
rect 521010 347052 521016 347064
rect 516192 347024 521016 347052
rect 516192 347012 516198 347024
rect 521010 347012 521016 347024
rect 521068 347012 521074 347064
rect 444374 346672 444380 346724
rect 444432 346712 444438 346724
rect 446398 346712 446404 346724
rect 444432 346684 446404 346712
rect 444432 346672 444438 346684
rect 446398 346672 446404 346684
rect 446456 346672 446462 346724
rect 445110 346604 445116 346656
rect 445168 346644 445174 346656
rect 446214 346644 446220 346656
rect 445168 346616 446220 346644
rect 445168 346604 445174 346616
rect 446214 346604 446220 346616
rect 446272 346604 446278 346656
rect 516226 346332 516232 346384
rect 516284 346372 516290 346384
rect 523218 346372 523224 346384
rect 516284 346344 523224 346372
rect 516284 346332 516290 346344
rect 523218 346332 523224 346344
rect 523276 346332 523282 346384
rect 370958 346264 370964 346316
rect 371016 346304 371022 346316
rect 374454 346304 374460 346316
rect 371016 346276 374460 346304
rect 371016 346264 371022 346276
rect 374454 346264 374460 346276
rect 374512 346264 374518 346316
rect 516134 346264 516140 346316
rect 516192 346304 516198 346316
rect 519538 346304 519544 346316
rect 516192 346276 519544 346304
rect 516192 346264 516198 346276
rect 519538 346264 519544 346276
rect 519596 346304 519602 346316
rect 522022 346304 522028 346316
rect 519596 346276 522028 346304
rect 519596 346264 519602 346276
rect 522022 346264 522028 346276
rect 522080 346264 522086 346316
rect 370222 345176 370228 345228
rect 370280 345216 370286 345228
rect 373074 345216 373080 345228
rect 370280 345188 373080 345216
rect 370280 345176 370286 345188
rect 373074 345176 373080 345188
rect 373132 345176 373138 345228
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 277486 345080 277492 345092
rect 3384 345052 277492 345080
rect 3384 345040 3390 345052
rect 277486 345040 277492 345052
rect 277544 345040 277550 345092
rect 516134 344292 516140 344344
rect 516192 344332 516198 344344
rect 519630 344332 519636 344344
rect 516192 344304 519636 344332
rect 516192 344292 516198 344304
rect 519630 344292 519636 344304
rect 519688 344332 519694 344344
rect 521838 344332 521844 344344
rect 519688 344304 521844 344332
rect 519688 344292 519694 344304
rect 521838 344292 521844 344304
rect 521896 344292 521902 344344
rect 445478 344156 445484 344208
rect 445536 344196 445542 344208
rect 447318 344196 447324 344208
rect 445536 344168 447324 344196
rect 445536 344156 445542 344168
rect 447318 344156 447324 344168
rect 447376 344156 447382 344208
rect 370958 343952 370964 344004
rect 371016 343992 371022 344004
rect 375650 343992 375656 344004
rect 371016 343964 375656 343992
rect 371016 343952 371022 343964
rect 375650 343952 375656 343964
rect 375708 343952 375714 344004
rect 444374 343884 444380 343936
rect 444432 343924 444438 343936
rect 449342 343924 449348 343936
rect 444432 343896 449348 343924
rect 444432 343884 444438 343896
rect 449342 343884 449348 343896
rect 449400 343884 449406 343936
rect 514754 343544 514760 343596
rect 514812 343584 514818 343596
rect 524690 343584 524696 343596
rect 514812 343556 524696 343584
rect 514812 343544 514818 343556
rect 524690 343544 524696 343556
rect 524748 343544 524754 343596
rect 370958 342864 370964 342916
rect 371016 342904 371022 342916
rect 372706 342904 372712 342916
rect 371016 342876 372712 342904
rect 371016 342864 371022 342876
rect 372706 342864 372712 342876
rect 372764 342904 372770 342916
rect 377306 342904 377312 342916
rect 372764 342876 377312 342904
rect 372764 342864 372770 342876
rect 377306 342864 377312 342876
rect 377364 342864 377370 342916
rect 443638 342252 443644 342304
rect 443696 342292 443702 342304
rect 444650 342292 444656 342304
rect 443696 342264 444656 342292
rect 443696 342252 443702 342264
rect 444650 342252 444656 342264
rect 444708 342252 444714 342304
rect 445110 342252 445116 342304
rect 445168 342292 445174 342304
rect 447042 342292 447048 342304
rect 445168 342264 447048 342292
rect 445168 342252 445174 342264
rect 447042 342252 447048 342264
rect 447100 342252 447106 342304
rect 447594 342184 447600 342236
rect 447652 342224 447658 342236
rect 447652 342196 451274 342224
rect 447652 342184 447658 342196
rect 451246 342088 451274 342196
rect 514754 342088 514760 342100
rect 451246 342060 514760 342088
rect 514754 342048 514760 342060
rect 514812 342048 514818 342100
rect 516134 341708 516140 341760
rect 516192 341748 516198 341760
rect 520366 341748 520372 341760
rect 516192 341720 520372 341748
rect 516192 341708 516198 341720
rect 520366 341708 520372 341720
rect 520424 341708 520430 341760
rect 441614 340892 441620 340944
rect 441672 340932 441678 340944
rect 447594 340932 447600 340944
rect 441672 340904 447600 340932
rect 441672 340892 441678 340904
rect 447594 340892 447600 340904
rect 447652 340892 447658 340944
rect 446398 340824 446404 340876
rect 446456 340864 446462 340876
rect 516410 340864 516416 340876
rect 446456 340836 516416 340864
rect 446456 340824 446462 340836
rect 516410 340824 516416 340836
rect 516468 340824 516474 340876
rect 472618 340756 472624 340808
rect 472676 340796 472682 340808
rect 513374 340796 513380 340808
rect 472676 340768 513380 340796
rect 472676 340756 472682 340768
rect 513374 340756 513380 340768
rect 513432 340756 513438 340808
rect 445478 340552 445484 340604
rect 445536 340592 445542 340604
rect 447226 340592 447232 340604
rect 445536 340564 447232 340592
rect 445536 340552 445542 340564
rect 447226 340552 447232 340564
rect 447284 340552 447290 340604
rect 444558 339464 444564 339516
rect 444616 339504 444622 339516
rect 471238 339504 471244 339516
rect 444616 339476 471244 339504
rect 444616 339464 444622 339476
rect 471238 339464 471244 339476
rect 471296 339504 471302 339516
rect 472618 339504 472624 339516
rect 471296 339476 472624 339504
rect 471296 339464 471302 339476
rect 472618 339464 472624 339476
rect 472676 339464 472682 339516
rect 368934 339192 368940 339244
rect 368992 339232 368998 339244
rect 369302 339232 369308 339244
rect 368992 339204 369308 339232
rect 368992 339192 368998 339204
rect 369302 339192 369308 339204
rect 369360 339192 369366 339244
rect 506842 338036 506848 338088
rect 506900 338076 506906 338088
rect 507762 338076 507768 338088
rect 506900 338048 507768 338076
rect 506900 338036 506906 338048
rect 507762 338036 507768 338048
rect 507820 338076 507826 338088
rect 513466 338076 513472 338088
rect 507820 338048 513472 338076
rect 507820 338036 507826 338048
rect 513466 338036 513472 338048
rect 513524 338036 513530 338088
rect 512914 337696 512920 337748
rect 512972 337736 512978 337748
rect 514754 337736 514760 337748
rect 512972 337708 514760 337736
rect 512972 337696 512978 337708
rect 514754 337696 514760 337708
rect 514812 337696 514818 337748
rect 322198 337424 322204 337476
rect 322256 337464 322262 337476
rect 366910 337464 366916 337476
rect 322256 337436 366916 337464
rect 322256 337424 322262 337436
rect 366910 337424 366916 337436
rect 366968 337424 366974 337476
rect 431218 337424 431224 337476
rect 431276 337464 431282 337476
rect 438946 337464 438952 337476
rect 431276 337436 438952 337464
rect 431276 337424 431282 337436
rect 438946 337424 438952 337436
rect 439004 337424 439010 337476
rect 300762 337356 300768 337408
rect 300820 337396 300826 337408
rect 510890 337396 510896 337408
rect 300820 337368 510896 337396
rect 300820 337356 300826 337368
rect 510890 337356 510896 337368
rect 510948 337356 510954 337408
rect 246942 330488 246948 330540
rect 247000 330528 247006 330540
rect 331214 330528 331220 330540
rect 247000 330500 331220 330528
rect 247000 330488 247006 330500
rect 331214 330488 331220 330500
rect 331272 330488 331278 330540
rect 41322 327700 41328 327752
rect 41380 327740 41386 327752
rect 258074 327740 258080 327752
rect 41380 327712 258080 327740
rect 41380 327700 41386 327712
rect 258074 327700 258080 327712
rect 258132 327700 258138 327752
rect 523034 326380 523040 326392
rect 451246 326352 523040 326380
rect 443638 326272 443644 326324
rect 443696 326312 443702 326324
rect 444190 326312 444196 326324
rect 443696 326284 444196 326312
rect 443696 326272 443702 326284
rect 444190 326272 444196 326284
rect 444248 326312 444254 326324
rect 451246 326312 451274 326352
rect 523034 326340 523040 326352
rect 523092 326340 523098 326392
rect 444248 326284 451274 326312
rect 444248 326272 444254 326284
rect 219342 324300 219348 324352
rect 219400 324340 219406 324352
rect 579614 324340 579620 324352
rect 219400 324312 579620 324340
rect 219400 324300 219406 324312
rect 579614 324300 579620 324312
rect 579672 324300 579678 324352
rect 378042 322192 378048 322244
rect 378100 322232 378106 322244
rect 525886 322232 525892 322244
rect 378100 322204 525892 322232
rect 378100 322192 378106 322204
rect 525886 322192 525892 322204
rect 525944 322192 525950 322244
rect 377398 321580 377404 321632
rect 377456 321620 377462 321632
rect 378042 321620 378048 321632
rect 377456 321592 378048 321620
rect 377456 321580 377462 321592
rect 378042 321580 378048 321592
rect 378100 321580 378106 321632
rect 373350 318860 373356 318912
rect 373408 318900 373414 318912
rect 373810 318900 373816 318912
rect 373408 318872 373816 318900
rect 373408 318860 373414 318872
rect 373810 318860 373816 318872
rect 373868 318900 373874 318912
rect 373868 318872 373994 318900
rect 373868 318860 373874 318872
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 278774 318832 278780 318844
rect 3476 318804 278780 318832
rect 3476 318792 3482 318804
rect 278774 318792 278780 318804
rect 278832 318792 278838 318844
rect 373966 318832 373994 318872
rect 441982 318832 441988 318844
rect 373966 318804 441988 318832
rect 441982 318792 441988 318804
rect 442040 318832 442046 318844
rect 443270 318832 443276 318844
rect 442040 318804 443276 318832
rect 442040 318792 442046 318804
rect 443270 318792 443276 318804
rect 443328 318792 443334 318844
rect 395338 318724 395344 318776
rect 395396 318764 395402 318776
rect 395982 318764 395988 318776
rect 395396 318736 395988 318764
rect 395396 318724 395402 318736
rect 395982 318724 395988 318736
rect 396040 318724 396046 318776
rect 395338 318044 395344 318096
rect 395396 318084 395402 318096
rect 521654 318084 521660 318096
rect 395396 318056 521660 318084
rect 395396 318044 395402 318056
rect 521654 318044 521660 318056
rect 521712 318044 521718 318096
rect 379422 315256 379428 315308
rect 379480 315296 379486 315308
rect 524506 315296 524512 315308
rect 379480 315268 524512 315296
rect 379480 315256 379486 315268
rect 524506 315256 524512 315268
rect 524564 315256 524570 315308
rect 378778 314644 378784 314696
rect 378836 314684 378842 314696
rect 379422 314684 379428 314696
rect 378836 314656 379428 314684
rect 378836 314644 378842 314656
rect 379422 314644 379428 314656
rect 379480 314644 379486 314696
rect 373258 313896 373264 313948
rect 373316 313936 373322 313948
rect 446214 313936 446220 313948
rect 373316 313908 446220 313936
rect 373316 313896 373322 313908
rect 446214 313896 446220 313908
rect 446272 313896 446278 313948
rect 220630 311856 220636 311908
rect 220688 311896 220694 311908
rect 580166 311896 580172 311908
rect 220688 311868 580172 311896
rect 220688 311856 220694 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 385770 310088 385776 310140
rect 385828 310128 385834 310140
rect 386322 310128 386328 310140
rect 385828 310100 386328 310128
rect 385828 310088 385834 310100
rect 386322 310088 386328 310100
rect 386380 310088 386386 310140
rect 386322 309748 386328 309800
rect 386380 309788 386386 309800
rect 527174 309788 527180 309800
rect 386380 309760 527180 309788
rect 386380 309748 386386 309760
rect 527174 309748 527180 309760
rect 527232 309748 527238 309800
rect 376018 309068 376024 309120
rect 376076 309108 376082 309120
rect 441890 309108 441896 309120
rect 376076 309080 441896 309108
rect 376076 309068 376082 309080
rect 441890 309068 441896 309080
rect 441948 309108 441954 309120
rect 444558 309108 444564 309120
rect 441948 309080 444564 309108
rect 441948 309068 441954 309080
rect 444558 309068 444564 309080
rect 444616 309068 444622 309120
rect 244458 307164 244464 307216
rect 244516 307204 244522 307216
rect 396718 307204 396724 307216
rect 244516 307176 396724 307204
rect 244516 307164 244522 307176
rect 396718 307164 396724 307176
rect 396776 307164 396782 307216
rect 241882 307096 241888 307148
rect 241940 307136 241946 307148
rect 461578 307136 461584 307148
rect 241940 307108 461584 307136
rect 241940 307096 241946 307108
rect 461578 307096 461584 307108
rect 461636 307096 461642 307148
rect 239306 307028 239312 307080
rect 239364 307068 239370 307080
rect 526438 307068 526444 307080
rect 239364 307040 526444 307068
rect 239364 307028 239370 307040
rect 526438 307028 526444 307040
rect 526496 307028 526502 307080
rect 248690 306008 248696 306060
rect 248748 306048 248754 306060
rect 295978 306048 295984 306060
rect 248748 306020 295984 306048
rect 248748 306008 248754 306020
rect 295978 306008 295984 306020
rect 296036 306008 296042 306060
rect 171042 305940 171048 305992
rect 171100 305980 171106 305992
rect 253750 305980 253756 305992
rect 171100 305952 253756 305980
rect 171100 305940 171106 305952
rect 253750 305940 253756 305952
rect 253808 305940 253814 305992
rect 246114 305872 246120 305924
rect 246172 305912 246178 305924
rect 359458 305912 359464 305924
rect 246172 305884 359464 305912
rect 246172 305872 246178 305884
rect 359458 305872 359464 305884
rect 359516 305872 359522 305924
rect 106182 305804 106188 305856
rect 106240 305844 106246 305856
rect 256234 305844 256240 305856
rect 106240 305816 256240 305844
rect 106240 305804 106246 305816
rect 256234 305804 256240 305816
rect 256292 305804 256298 305856
rect 243538 305736 243544 305788
rect 243596 305776 243602 305788
rect 429194 305776 429200 305788
rect 243596 305748 429200 305776
rect 243596 305736 243602 305748
rect 429194 305736 429200 305748
rect 429252 305736 429258 305788
rect 228266 305668 228272 305720
rect 228324 305708 228330 305720
rect 582374 305708 582380 305720
rect 228324 305680 582380 305708
rect 228324 305668 228330 305680
rect 582374 305668 582380 305680
rect 582432 305668 582438 305720
rect 226610 305600 226616 305652
rect 226668 305640 226674 305652
rect 582466 305640 582472 305652
rect 226668 305612 582472 305640
rect 226668 305600 226674 305612
rect 582466 305600 582472 305612
rect 582524 305600 582530 305652
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 280890 305028 280896 305040
rect 3292 305000 280896 305028
rect 3292 304988 3298 305000
rect 280890 304988 280896 305000
rect 280948 304988 280954 305040
rect 233142 304784 233148 304836
rect 233200 304824 233206 304836
rect 251174 304824 251180 304836
rect 233200 304796 251180 304824
rect 233200 304784 233206 304796
rect 251174 304784 251180 304796
rect 251232 304784 251238 304836
rect 241054 304716 241060 304768
rect 241112 304756 241118 304768
rect 494054 304756 494060 304768
rect 241112 304728 494060 304756
rect 241112 304716 241118 304728
rect 494054 304716 494060 304728
rect 494112 304716 494118 304768
rect 238478 304648 238484 304700
rect 238536 304688 238542 304700
rect 558914 304688 558920 304700
rect 238536 304660 558920 304688
rect 238536 304648 238542 304660
rect 558914 304648 558920 304660
rect 558972 304648 558978 304700
rect 232590 304580 232596 304632
rect 232648 304620 232654 304632
rect 580258 304620 580264 304632
rect 232648 304592 580264 304620
rect 232648 304580 232654 304592
rect 580258 304580 580264 304592
rect 580316 304580 580322 304632
rect 230842 304512 230848 304564
rect 230900 304552 230906 304564
rect 580350 304552 580356 304564
rect 230900 304524 580356 304552
rect 230900 304512 230906 304524
rect 580350 304512 580356 304524
rect 580408 304512 580414 304564
rect 224954 304444 224960 304496
rect 225012 304484 225018 304496
rect 580534 304484 580540 304496
rect 225012 304456 580540 304484
rect 225012 304444 225018 304456
rect 580534 304444 580540 304456
rect 580592 304444 580598 304496
rect 224034 304376 224040 304428
rect 224092 304416 224098 304428
rect 580442 304416 580448 304428
rect 224092 304388 580448 304416
rect 224092 304376 224098 304388
rect 580442 304376 580448 304388
rect 580500 304376 580506 304428
rect 222378 304308 222384 304360
rect 222436 304348 222442 304360
rect 580626 304348 580632 304360
rect 222436 304320 580632 304348
rect 222436 304308 222442 304320
rect 580626 304308 580632 304320
rect 580684 304308 580690 304360
rect 220722 304240 220728 304292
rect 220780 304280 220786 304292
rect 580718 304280 580724 304292
rect 220780 304252 580724 304280
rect 220780 304240 220786 304252
rect 580718 304240 580724 304252
rect 580776 304240 580782 304292
rect 262214 303220 262220 303272
rect 262272 303260 262278 303272
rect 262766 303260 262772 303272
rect 262272 303232 262772 303260
rect 262272 303220 262278 303232
rect 262766 303220 262772 303232
rect 262824 303220 262830 303272
rect 274634 303220 274640 303272
rect 274692 303260 274698 303272
rect 275462 303260 275468 303272
rect 274692 303232 275468 303260
rect 274692 303220 274698 303232
rect 275462 303220 275468 303232
rect 275520 303220 275526 303272
rect 277394 303220 277400 303272
rect 277452 303260 277458 303272
rect 278038 303260 278044 303272
rect 277452 303232 278044 303260
rect 277452 303220 277458 303232
rect 278038 303220 278044 303232
rect 278096 303220 278102 303272
rect 212166 303152 212172 303204
rect 212224 303192 212230 303204
rect 536098 303192 536104 303204
rect 212224 303164 536104 303192
rect 212224 303152 212230 303164
rect 536098 303152 536104 303164
rect 536156 303152 536162 303204
rect 207106 303084 207112 303136
rect 207164 303124 207170 303136
rect 533338 303124 533344 303136
rect 207164 303096 533344 303124
rect 207164 303084 207170 303096
rect 533338 303084 533344 303096
rect 533396 303084 533402 303136
rect 204622 303016 204628 303068
rect 204680 303056 204686 303068
rect 530578 303056 530584 303068
rect 204680 303028 530584 303056
rect 204680 303016 204686 303028
rect 530578 303016 530584 303028
rect 530636 303016 530642 303068
rect 43438 302948 43444 303000
rect 43496 302988 43502 303000
rect 296070 302988 296076 303000
rect 43496 302960 296076 302988
rect 43496 302948 43502 302960
rect 296070 302948 296076 302960
rect 296128 302948 296134 303000
rect 28258 302880 28264 302932
rect 28316 302920 28322 302932
rect 285950 302920 285956 302932
rect 28316 302892 285956 302920
rect 28316 302880 28322 302892
rect 285950 302880 285956 302892
rect 286008 302880 286014 302932
rect 29638 302812 29644 302864
rect 29696 302852 29702 302864
rect 288526 302852 288532 302864
rect 29696 302824 288532 302852
rect 29696 302812 29702 302824
rect 288526 302812 288532 302824
rect 288584 302812 288590 302864
rect 299474 302812 299480 302864
rect 299532 302852 299538 302864
rect 300762 302852 300768 302864
rect 299532 302824 300768 302852
rect 299532 302812 299538 302824
rect 300762 302812 300768 302824
rect 300820 302812 300826 302864
rect 32398 302744 32404 302796
rect 32456 302784 32462 302796
rect 293586 302784 293592 302796
rect 32456 302756 293592 302784
rect 32456 302744 32462 302756
rect 293586 302744 293592 302756
rect 293644 302744 293650 302796
rect 26878 302676 26884 302728
rect 26936 302716 26942 302728
rect 295242 302716 295248 302728
rect 26936 302688 295248 302716
rect 26936 302676 26942 302688
rect 295242 302676 295248 302688
rect 295300 302676 295306 302728
rect 4798 302608 4804 302660
rect 4856 302648 4862 302660
rect 291010 302648 291016 302660
rect 4856 302620 291016 302648
rect 4856 302608 4862 302620
rect 291010 302608 291016 302620
rect 291068 302608 291074 302660
rect 211338 302540 211344 302592
rect 211396 302580 211402 302592
rect 522298 302580 522304 302592
rect 211396 302552 522304 302580
rect 211396 302540 211402 302552
rect 522298 302540 522304 302552
rect 522356 302540 522362 302592
rect 208854 302472 208860 302524
rect 208912 302512 208918 302524
rect 520918 302512 520924 302524
rect 208912 302484 520924 302512
rect 208912 302472 208918 302484
rect 520918 302472 520924 302484
rect 520976 302472 520982 302524
rect 202046 302404 202052 302456
rect 202104 302444 202110 302456
rect 525058 302444 525064 302456
rect 202104 302416 525064 302444
rect 202104 302404 202110 302416
rect 525058 302404 525064 302416
rect 525116 302404 525122 302456
rect 296990 302336 296996 302388
rect 297048 302376 297054 302388
rect 297048 302348 306374 302376
rect 297048 302336 297054 302348
rect 297818 302268 297824 302320
rect 297876 302308 297882 302320
rect 306346 302308 306374 302348
rect 307018 302308 307024 302320
rect 297876 302280 305776 302308
rect 306346 302280 307024 302308
rect 297876 302268 297882 302280
rect 298646 302200 298652 302252
rect 298704 302240 298710 302252
rect 305638 302240 305644 302252
rect 298704 302212 305644 302240
rect 298704 302200 298710 302212
rect 305638 302200 305644 302212
rect 305696 302200 305702 302252
rect 305748 302240 305776 302280
rect 307018 302268 307024 302280
rect 307076 302268 307082 302320
rect 309778 302240 309784 302252
rect 305748 302212 309784 302240
rect 309778 302200 309784 302212
rect 309836 302200 309842 302252
rect 229186 302064 229192 302116
rect 229244 302104 229250 302116
rect 230382 302104 230388 302116
rect 229244 302076 230388 302104
rect 229244 302064 229250 302076
rect 230382 302064 230388 302076
rect 230440 302064 230446 302116
rect 199378 301588 199384 301640
rect 199436 301628 199442 301640
rect 284202 301628 284208 301640
rect 199436 301600 284208 301628
rect 199436 301588 199442 301600
rect 284202 301588 284208 301600
rect 284260 301588 284266 301640
rect 210510 301520 210516 301572
rect 210568 301560 210574 301572
rect 301498 301560 301504 301572
rect 210568 301532 301504 301560
rect 210568 301520 210574 301532
rect 301498 301520 301504 301532
rect 301556 301520 301562 301572
rect 215570 301452 215576 301504
rect 215628 301492 215634 301504
rect 312538 301492 312544 301504
rect 215628 301464 312544 301492
rect 215628 301452 215634 301464
rect 312538 301452 312544 301464
rect 312596 301452 312602 301504
rect 206278 301384 206284 301436
rect 206336 301424 206342 301436
rect 318058 301424 318064 301436
rect 206336 301396 318064 301424
rect 206336 301384 206342 301396
rect 318058 301384 318064 301396
rect 318116 301384 318122 301436
rect 201218 301316 201224 301368
rect 201276 301356 201282 301368
rect 313918 301356 313924 301368
rect 201276 301328 313924 301356
rect 201276 301316 201282 301328
rect 313918 301316 313924 301328
rect 313976 301316 313982 301368
rect 152458 301248 152464 301300
rect 152516 301288 152522 301300
rect 287606 301288 287612 301300
rect 152516 301260 287612 301288
rect 152516 301248 152522 301260
rect 287606 301248 287612 301260
rect 287664 301248 287670 301300
rect 156598 301180 156604 301232
rect 156656 301220 156662 301232
rect 294414 301220 294420 301232
rect 156656 301192 294420 301220
rect 156656 301180 156662 301192
rect 294414 301180 294420 301192
rect 294472 301180 294478 301232
rect 148318 301112 148324 301164
rect 148376 301152 148382 301164
rect 292758 301152 292764 301164
rect 148376 301124 292764 301152
rect 148376 301112 148382 301124
rect 292758 301112 292764 301124
rect 292816 301112 292822 301164
rect 10318 301044 10324 301096
rect 10376 301084 10382 301096
rect 281718 301084 281724 301096
rect 10376 301056 281724 301084
rect 10376 301044 10382 301056
rect 281718 301044 281724 301056
rect 281776 301044 281782 301096
rect 214742 300976 214748 301028
rect 214800 301016 214806 301028
rect 519538 301016 519544 301028
rect 214800 300988 519544 301016
rect 214800 300976 214806 300988
rect 519538 300976 519544 300988
rect 519596 300976 519602 301028
rect 202874 300908 202880 300960
rect 202932 300948 202938 300960
rect 582466 300948 582472 300960
rect 202932 300920 582472 300948
rect 202932 300908 202938 300920
rect 582466 300908 582472 300920
rect 582524 300908 582530 300960
rect 200390 300840 200396 300892
rect 200448 300880 200454 300892
rect 582374 300880 582380 300892
rect 200448 300852 582380 300880
rect 200448 300840 200454 300852
rect 582374 300840 582380 300852
rect 582432 300840 582438 300892
rect 219802 300228 219808 300280
rect 219860 300268 219866 300280
rect 220630 300268 220636 300280
rect 219860 300240 220636 300268
rect 219860 300228 219866 300240
rect 220630 300228 220636 300240
rect 220688 300228 220694 300280
rect 233418 300228 233424 300280
rect 233476 300268 233482 300280
rect 234430 300268 234436 300280
rect 233476 300240 234436 300268
rect 233476 300228 233482 300240
rect 234430 300228 234436 300240
rect 234488 300228 234494 300280
rect 237650 300228 237656 300280
rect 237708 300268 237714 300280
rect 238570 300268 238576 300280
rect 237708 300240 238576 300268
rect 237708 300228 237714 300240
rect 238570 300228 238576 300240
rect 238628 300228 238634 300280
rect 240134 300228 240140 300280
rect 240192 300268 240198 300280
rect 241330 300268 241336 300280
rect 240192 300240 241336 300268
rect 240192 300228 240198 300240
rect 241330 300228 241336 300240
rect 241388 300228 241394 300280
rect 205450 300160 205456 300212
rect 205508 300200 205514 300212
rect 311158 300200 311164 300212
rect 205508 300172 311164 300200
rect 205508 300160 205514 300172
rect 311158 300160 311164 300172
rect 311216 300160 311222 300212
rect 203702 300092 203708 300144
rect 203760 300132 203766 300144
rect 316678 300132 316684 300144
rect 203760 300104 316684 300132
rect 203760 300092 203766 300104
rect 316678 300092 316684 300104
rect 316736 300092 316742 300144
rect 155218 300024 155224 300076
rect 155276 300064 155282 300076
rect 284846 300064 284852 300076
rect 155276 300036 284852 300064
rect 155276 300024 155282 300036
rect 284846 300024 284852 300036
rect 284904 300024 284910 300076
rect 159358 299956 159364 300008
rect 159416 299996 159422 300008
rect 289078 299996 289084 300008
rect 159416 299968 289084 299996
rect 159416 299956 159422 299968
rect 289078 299956 289084 299968
rect 289136 299956 289142 300008
rect 157978 299888 157984 299940
rect 158036 299928 158042 299940
rect 291470 299928 291476 299940
rect 158036 299900 291476 299928
rect 158036 299888 158042 299900
rect 291470 299888 291476 299900
rect 291528 299888 291534 299940
rect 151078 299820 151084 299872
rect 151136 299860 151142 299872
rect 289814 299860 289820 299872
rect 151136 299832 289820 299860
rect 151136 299820 151142 299832
rect 289814 299820 289820 299832
rect 289872 299820 289878 299872
rect 371418 299820 371424 299872
rect 371476 299860 371482 299872
rect 375282 299860 375288 299872
rect 371476 299832 375288 299860
rect 371476 299820 371482 299832
rect 375282 299820 375288 299832
rect 375340 299820 375346 299872
rect 11698 299752 11704 299804
rect 11756 299792 11762 299804
rect 286502 299792 286508 299804
rect 11756 299764 286508 299792
rect 11756 299752 11762 299764
rect 286502 299752 286508 299764
rect 286560 299752 286566 299804
rect 213362 299684 213368 299736
rect 213420 299724 213426 299736
rect 515398 299724 515404 299736
rect 213420 299696 515404 299724
rect 213420 299684 213426 299696
rect 515398 299684 515404 299696
rect 515456 299684 515462 299736
rect 210050 299616 210056 299668
rect 210108 299656 210114 299668
rect 518158 299656 518164 299668
rect 210108 299628 518164 299656
rect 210108 299616 210114 299628
rect 518158 299616 518164 299628
rect 518216 299616 518222 299668
rect 208210 299548 208216 299600
rect 208268 299588 208274 299600
rect 526438 299588 526444 299600
rect 208268 299560 526444 299588
rect 208268 299548 208274 299560
rect 526438 299548 526444 299560
rect 526496 299548 526502 299600
rect 218514 299480 218520 299532
rect 218572 299520 218578 299532
rect 580166 299520 580172 299532
rect 218572 299492 580172 299520
rect 218572 299480 218578 299492
rect 580166 299480 580172 299492
rect 580224 299480 580230 299532
rect 214006 299412 214012 299464
rect 214064 299452 214070 299464
rect 214064 299424 249794 299452
rect 214064 299412 214070 299424
rect 208366 299356 231854 299384
rect 208366 298840 208394 299356
rect 214006 299316 214012 299328
rect 205606 298812 208394 298840
rect 211126 299288 214012 299316
rect 205606 298772 205634 298812
rect 200086 298744 205634 298772
rect 198458 298528 198464 298580
rect 198516 298568 198522 298580
rect 200086 298568 200114 298744
rect 198516 298540 200114 298568
rect 198516 298528 198522 298540
rect 3878 298460 3884 298512
rect 3936 298500 3942 298512
rect 211126 298500 211154 299288
rect 214006 299276 214012 299288
rect 214064 299276 214070 299328
rect 214558 299276 214564 299328
rect 214616 299276 214622 299328
rect 214650 299276 214656 299328
rect 214708 299276 214714 299328
rect 216030 299276 216036 299328
rect 216088 299276 216094 299328
rect 216858 299276 216864 299328
rect 216916 299276 216922 299328
rect 216950 299276 216956 299328
rect 217008 299276 217014 299328
rect 217594 299276 217600 299328
rect 217652 299316 217658 299328
rect 217652 299288 224264 299316
rect 217652 299276 217658 299288
rect 3936 298472 211154 298500
rect 3936 298460 3942 298472
rect 3418 298392 3424 298444
rect 3476 298432 3482 298444
rect 214576 298432 214604 299276
rect 3476 298404 204254 298432
rect 3476 298392 3482 298404
rect 3510 298324 3516 298376
rect 3568 298364 3574 298376
rect 3568 298336 200114 298364
rect 3568 298324 3574 298336
rect 200086 298228 200114 298336
rect 204226 298296 204254 298404
rect 211126 298404 214604 298432
rect 211126 298296 211154 298404
rect 204226 298268 211154 298296
rect 200086 298200 204254 298228
rect 204226 298024 204254 298200
rect 204226 297996 209774 298024
rect 209746 297820 209774 297996
rect 214668 297820 214696 299276
rect 209746 297792 214696 297820
rect 216048 297616 216076 299276
rect 216876 298500 216904 299276
rect 216968 299248 216996 299276
rect 216968 299220 220124 299248
rect 220096 298568 220124 299220
rect 224236 298908 224264 299288
rect 224402 299276 224408 299328
rect 224460 299316 224466 299328
rect 224460 299288 230474 299316
rect 224460 299276 224466 299288
rect 224236 298880 224954 298908
rect 224926 298636 224954 298880
rect 230446 298704 230474 299288
rect 231826 299044 231854 299356
rect 231826 299016 238754 299044
rect 238726 298908 238754 299016
rect 238726 298880 247724 298908
rect 238726 298812 247632 298840
rect 238726 298704 238754 298812
rect 230446 298676 238754 298704
rect 247604 298636 247632 298812
rect 247696 298704 247724 298880
rect 249766 298840 249794 299424
rect 282638 299412 282644 299464
rect 282696 299452 282702 299464
rect 283466 299452 283472 299464
rect 282696 299424 283472 299452
rect 282696 299412 282702 299424
rect 283466 299412 283472 299424
rect 283524 299412 283530 299464
rect 280172 299356 285674 299384
rect 279694 299316 279700 299328
rect 277366 299288 279700 299316
rect 259426 299084 269114 299112
rect 259426 298976 259454 299084
rect 259656 299016 268056 299044
rect 259656 298976 259684 299016
rect 258046 298948 259454 298976
rect 259564 298948 259684 298976
rect 258046 298840 258074 298948
rect 259564 298908 259592 298948
rect 268028 298908 268056 299016
rect 269086 298976 269114 299084
rect 277366 298976 277394 299288
rect 279694 299276 279700 299288
rect 279752 299276 279758 299328
rect 280172 299112 280200 299356
rect 282270 299276 282276 299328
rect 282328 299276 282334 299328
rect 282638 299276 282644 299328
rect 282696 299276 282702 299328
rect 283006 299276 283012 299328
rect 283064 299276 283070 299328
rect 283466 299276 283472 299328
rect 283524 299316 283530 299328
rect 283524 299288 284294 299316
rect 283524 299276 283530 299288
rect 269086 298948 277394 298976
rect 278608 299084 280200 299112
rect 278608 298908 278636 299084
rect 282288 299044 282316 299276
rect 259472 298880 259592 298908
rect 259748 298880 267872 298908
rect 268028 298880 278636 298908
rect 279252 299016 282316 299044
rect 259472 298840 259500 298880
rect 249766 298812 258074 298840
rect 258276 298812 259500 298840
rect 249766 298744 258074 298772
rect 249766 298704 249794 298744
rect 247696 298676 249794 298704
rect 258046 298636 258074 298744
rect 258276 298636 258304 298812
rect 259748 298772 259776 298880
rect 267844 298840 267872 298880
rect 259426 298744 259776 298772
rect 261220 298812 264376 298840
rect 267844 298812 276060 298840
rect 259426 298704 259454 298744
rect 224926 298608 230474 298636
rect 247604 298608 249794 298636
rect 258046 298608 258304 298636
rect 258368 298676 259454 298704
rect 220096 298540 227714 298568
rect 216876 298472 226334 298500
rect 226306 297888 226334 298472
rect 227686 298092 227714 298540
rect 230446 298296 230474 298608
rect 249766 298568 249794 298608
rect 258368 298568 258396 298676
rect 231826 298540 242894 298568
rect 249766 298540 258396 298568
rect 231826 298296 231854 298540
rect 242866 298500 242894 298540
rect 242866 298472 249794 298500
rect 249766 298364 249794 298472
rect 261220 298364 261248 298812
rect 264348 298568 264376 298812
rect 276032 298772 276060 298812
rect 279252 298772 279280 299016
rect 264946 298744 274634 298772
rect 276032 298744 279280 298772
rect 264946 298568 264974 298744
rect 274606 298704 274634 298744
rect 282656 298704 282684 299276
rect 274606 298676 282684 298704
rect 264348 298540 264974 298568
rect 249766 298336 261248 298364
rect 262232 298472 262444 298500
rect 262232 298296 262260 298472
rect 262416 298432 262444 298472
rect 283024 298432 283052 299276
rect 262416 298404 262536 298432
rect 230446 298268 231854 298296
rect 240106 298268 249472 298296
rect 240106 298160 240134 298268
rect 229066 298132 231854 298160
rect 229066 298092 229094 298132
rect 227686 298064 229094 298092
rect 231826 298092 231854 298132
rect 233206 298132 234614 298160
rect 233206 298092 233234 298132
rect 231826 298064 233234 298092
rect 234586 298092 234614 298132
rect 235966 298132 240134 298160
rect 246684 298200 249380 298228
rect 235966 298092 235994 298132
rect 234586 298064 235994 298092
rect 236012 297996 237374 298024
rect 236012 297956 236040 297996
rect 234586 297928 236040 297956
rect 237346 297956 237374 297996
rect 237346 297928 238754 297956
rect 226306 297860 227714 297888
rect 227686 297684 227714 297860
rect 234586 297684 234614 297928
rect 227686 297656 234614 297684
rect 238726 297684 238754 297928
rect 246684 297684 246712 298200
rect 238726 297656 246712 297684
rect 247006 298132 249288 298160
rect 247006 297616 247034 298132
rect 249260 297956 249288 298132
rect 249352 298024 249380 298200
rect 249444 298160 249472 298268
rect 262140 298268 262260 298296
rect 262508 298296 262536 298404
rect 274606 298404 283052 298432
rect 274606 298364 274634 298404
rect 264946 298336 274634 298364
rect 284266 298364 284294 299288
rect 285646 298908 285674 299356
rect 375926 299072 375932 299124
rect 375984 299112 375990 299124
rect 376662 299112 376668 299124
rect 375984 299084 376668 299112
rect 375984 299072 375990 299084
rect 376662 299072 376668 299084
rect 376720 299072 376726 299124
rect 285646 298880 287054 298908
rect 287026 298772 287054 298880
rect 382274 298800 382280 298852
rect 382332 298840 382338 298852
rect 394602 298840 394608 298852
rect 382332 298812 394608 298840
rect 382332 298800 382338 298812
rect 394602 298800 394608 298812
rect 394660 298840 394666 298852
rect 516778 298840 516784 298852
rect 394660 298812 516784 298840
rect 394660 298800 394666 298812
rect 516778 298800 516784 298812
rect 516836 298800 516842 298852
rect 287026 298744 288434 298772
rect 288406 298568 288434 298744
rect 379422 298732 379428 298784
rect 379480 298772 379486 298784
rect 383562 298772 383568 298784
rect 379480 298744 383568 298772
rect 379480 298732 379486 298744
rect 383562 298732 383568 298744
rect 383620 298772 383626 298784
rect 516594 298772 516600 298784
rect 383620 298744 516600 298772
rect 383620 298732 383626 298744
rect 516594 298732 516600 298744
rect 516652 298732 516658 298784
rect 429838 298568 429844 298580
rect 288406 298540 429844 298568
rect 429838 298528 429844 298540
rect 429896 298528 429902 298580
rect 507762 298460 507768 298512
rect 507820 298500 507826 298512
rect 514202 298500 514208 298512
rect 507820 298472 514208 298500
rect 507820 298460 507826 298472
rect 514202 298460 514208 298472
rect 514260 298460 514266 298512
rect 382182 298392 382188 298444
rect 382240 298432 382246 298444
rect 516686 298432 516692 298444
rect 382240 298404 516692 298432
rect 382240 298392 382246 298404
rect 516686 298392 516692 298404
rect 516744 298392 516750 298444
rect 284266 298336 289814 298364
rect 264946 298296 264974 298336
rect 262508 298268 264974 298296
rect 289786 298296 289814 298336
rect 375926 298324 375932 298376
rect 375984 298364 375990 298376
rect 516502 298364 516508 298376
rect 375984 298336 516508 298364
rect 375984 298324 375990 298336
rect 516502 298324 516508 298336
rect 516560 298324 516566 298376
rect 580350 298296 580356 298308
rect 289786 298268 580356 298296
rect 249444 298132 251174 298160
rect 251146 298092 251174 298132
rect 262140 298092 262168 298268
rect 580350 298256 580356 298268
rect 580408 298256 580414 298308
rect 580442 298228 580448 298240
rect 251146 298064 262168 298092
rect 263888 298200 267872 298228
rect 249352 297996 262444 298024
rect 262416 297956 262444 297996
rect 263888 297956 263916 298200
rect 267844 298160 267872 298200
rect 271616 298200 280292 298228
rect 271616 298160 271644 298200
rect 280264 298160 280292 298200
rect 280540 298200 580448 298228
rect 280540 298160 280568 298200
rect 580442 298188 580448 298200
rect 580500 298188 580506 298240
rect 580258 298160 580264 298172
rect 267844 298132 268056 298160
rect 268028 298092 268056 298132
rect 268396 298132 271644 298160
rect 277366 298132 280154 298160
rect 280264 298132 280568 298160
rect 284956 298132 580264 298160
rect 268396 298092 268424 298132
rect 249260 297928 258074 297956
rect 262416 297928 263916 297956
rect 264946 298064 267872 298092
rect 268028 298064 268424 298092
rect 258046 297888 258074 297928
rect 264946 297888 264974 298064
rect 267844 297956 267872 298064
rect 258046 297860 264974 297888
rect 267752 297928 267872 297956
rect 267752 297820 267780 297928
rect 277366 297820 277394 298132
rect 280126 298024 280154 298132
rect 284956 298024 284984 298132
rect 580258 298120 580264 298132
rect 580316 298120 580322 298172
rect 441890 298052 441896 298104
rect 441948 298092 441954 298104
rect 442442 298092 442448 298104
rect 441948 298064 442448 298092
rect 441948 298052 441954 298064
rect 442442 298052 442448 298064
rect 442500 298052 442506 298104
rect 445294 298052 445300 298104
rect 445352 298092 445358 298104
rect 445662 298092 445668 298104
rect 445352 298064 445668 298092
rect 445352 298052 445358 298064
rect 445662 298052 445668 298064
rect 445720 298052 445726 298104
rect 280126 297996 284984 298024
rect 371326 297984 371332 298036
rect 371384 298024 371390 298036
rect 375190 298024 375196 298036
rect 371384 297996 375196 298024
rect 371384 297984 371390 297996
rect 375190 297984 375196 297996
rect 375248 297984 375254 298036
rect 445110 297984 445116 298036
rect 445168 298024 445174 298036
rect 445570 298024 445576 298036
rect 445168 297996 445576 298024
rect 445168 297984 445174 297996
rect 445570 297984 445576 297996
rect 445628 297984 445634 298036
rect 507854 297848 507860 297900
rect 507912 297888 507918 297900
rect 513742 297888 513748 297900
rect 507912 297860 513748 297888
rect 507912 297848 507918 297860
rect 513742 297848 513748 297860
rect 513800 297848 513806 297900
rect 267752 297792 277394 297820
rect 216048 297588 247034 297616
rect 442442 297576 442448 297628
rect 442500 297616 442506 297628
rect 442500 297588 451274 297616
rect 442500 297576 442506 297588
rect 444374 297508 444380 297560
rect 444432 297548 444438 297560
rect 446122 297548 446128 297560
rect 444432 297520 446128 297548
rect 444432 297508 444438 297520
rect 446122 297508 446128 297520
rect 446180 297508 446186 297560
rect 451246 297548 451274 297588
rect 516318 297548 516324 297560
rect 451246 297520 489914 297548
rect 303062 297440 303068 297492
rect 303120 297480 303126 297492
rect 369394 297480 369400 297492
rect 303120 297452 369400 297480
rect 303120 297440 303126 297452
rect 369394 297440 369400 297452
rect 369452 297440 369458 297492
rect 443270 297440 443276 297492
rect 443328 297480 443334 297492
rect 444282 297480 444288 297492
rect 443328 297452 444288 297480
rect 443328 297440 443334 297452
rect 444282 297440 444288 297452
rect 444340 297440 444346 297492
rect 489886 297480 489914 297520
rect 505066 297520 516324 297548
rect 505066 297480 505094 297520
rect 516318 297508 516324 297520
rect 516376 297508 516382 297560
rect 489886 297452 505094 297480
rect 302878 297372 302884 297424
rect 302936 297412 302942 297424
rect 369854 297412 369860 297424
rect 302936 297384 369860 297412
rect 302936 297372 302942 297384
rect 369854 297372 369860 297384
rect 369912 297372 369918 297424
rect 375190 297372 375196 297424
rect 375248 297412 375254 297424
rect 513374 297412 513380 297424
rect 375248 297384 513380 297412
rect 375248 297372 375254 297384
rect 513374 297372 513380 297384
rect 513432 297372 513438 297424
rect 448422 297304 448428 297356
rect 448480 297344 448486 297356
rect 517146 297344 517152 297356
rect 448480 297316 517152 297344
rect 448480 297304 448486 297316
rect 517146 297304 517152 297316
rect 517204 297304 517210 297356
rect 445386 297236 445392 297288
rect 445444 297276 445450 297288
rect 514110 297276 514116 297288
rect 445444 297248 514116 297276
rect 445444 297236 445450 297248
rect 514110 297236 514116 297248
rect 514168 297236 514174 297288
rect 445110 297168 445116 297220
rect 445168 297208 445174 297220
rect 513282 297208 513288 297220
rect 445168 297180 513288 297208
rect 445168 297168 445174 297180
rect 513282 297168 513288 297180
rect 513340 297168 513346 297220
rect 444926 297100 444932 297152
rect 444984 297140 444990 297152
rect 513926 297140 513932 297152
rect 444984 297112 513932 297140
rect 444984 297100 444990 297112
rect 513926 297100 513932 297112
rect 513984 297100 513990 297152
rect 444742 297032 444748 297084
rect 444800 297072 444806 297084
rect 513834 297072 513840 297084
rect 444800 297044 513840 297072
rect 444800 297032 444806 297044
rect 513834 297032 513840 297044
rect 513892 297032 513898 297084
rect 445662 296964 445668 297016
rect 445720 297004 445726 297016
rect 516410 297004 516416 297016
rect 445720 296976 516416 297004
rect 445720 296964 445726 296976
rect 516410 296964 516416 296976
rect 516468 296964 516474 297016
rect 444282 296896 444288 296948
rect 444340 296936 444346 296948
rect 516226 296936 516232 296948
rect 444340 296908 516232 296936
rect 444340 296896 444346 296908
rect 516226 296896 516232 296908
rect 516284 296896 516290 296948
rect 442258 296828 442264 296880
rect 442316 296868 442322 296880
rect 516134 296868 516140 296880
rect 442316 296840 516140 296868
rect 442316 296828 442322 296840
rect 516134 296828 516140 296840
rect 516192 296828 516198 296880
rect 371786 296760 371792 296812
rect 371844 296800 371850 296812
rect 371844 296772 373994 296800
rect 371844 296760 371850 296772
rect 373966 296732 373994 296772
rect 425698 296760 425704 296812
rect 425756 296800 425762 296812
rect 441706 296800 441712 296812
rect 425756 296772 441712 296800
rect 425756 296760 425762 296772
rect 441706 296760 441712 296772
rect 441764 296760 441770 296812
rect 375098 296732 375104 296744
rect 373966 296704 375104 296732
rect 375098 296692 375104 296704
rect 375156 296732 375162 296744
rect 513374 296732 513380 296744
rect 375156 296704 513380 296732
rect 375156 296692 375162 296704
rect 513374 296692 513380 296704
rect 513432 296692 513438 296744
rect 371234 296624 371240 296676
rect 371292 296664 371298 296676
rect 389082 296664 389088 296676
rect 371292 296636 389088 296664
rect 371292 296624 371298 296636
rect 389082 296624 389088 296636
rect 389140 296624 389146 296676
rect 390462 296556 390468 296608
rect 390520 296596 390526 296608
rect 513374 296596 513380 296608
rect 390520 296568 513380 296596
rect 390520 296556 390526 296568
rect 513374 296556 513380 296568
rect 513432 296596 513438 296608
rect 517238 296596 517244 296608
rect 513432 296568 517244 296596
rect 513432 296556 513438 296568
rect 517238 296556 517244 296568
rect 517296 296556 517302 296608
rect 378870 296488 378876 296540
rect 378928 296528 378934 296540
rect 443270 296528 443276 296540
rect 378928 296500 443276 296528
rect 378928 296488 378934 296500
rect 443270 296488 443276 296500
rect 443328 296488 443334 296540
rect 444374 296488 444380 296540
rect 444432 296528 444438 296540
rect 446030 296528 446036 296540
rect 444432 296500 446036 296528
rect 444432 296488 444438 296500
rect 446030 296488 446036 296500
rect 446088 296488 446094 296540
rect 389082 296420 389088 296472
rect 389140 296460 389146 296472
rect 513466 296460 513472 296472
rect 389140 296432 513472 296460
rect 389140 296420 389146 296432
rect 513466 296420 513472 296432
rect 513524 296420 513530 296472
rect 347682 296148 347688 296200
rect 347740 296188 347746 296200
rect 369394 296188 369400 296200
rect 347740 296160 369400 296188
rect 347740 296148 347746 296160
rect 369394 296148 369400 296160
rect 369452 296188 369458 296200
rect 371234 296188 371240 296200
rect 369452 296160 371240 296188
rect 369452 296148 369458 296160
rect 371234 296148 371240 296160
rect 371292 296148 371298 296200
rect 375282 296148 375288 296200
rect 375340 296188 375346 296200
rect 391934 296188 391940 296200
rect 375340 296160 391940 296188
rect 375340 296148 375346 296160
rect 391934 296148 391940 296160
rect 391992 296148 391998 296200
rect 372338 296080 372344 296132
rect 372396 296120 372402 296132
rect 390462 296120 390468 296132
rect 372396 296092 390468 296120
rect 372396 296080 372402 296092
rect 390462 296080 390468 296092
rect 390520 296080 390526 296132
rect 400674 296080 400680 296132
rect 400732 296120 400738 296132
rect 443638 296120 443644 296132
rect 400732 296092 443644 296120
rect 400732 296080 400738 296092
rect 443638 296080 443644 296092
rect 443696 296080 443702 296132
rect 358078 296012 358084 296064
rect 358136 296052 358142 296064
rect 371418 296052 371424 296064
rect 358136 296024 371424 296052
rect 358136 296012 358142 296024
rect 371418 296012 371424 296024
rect 371476 296012 371482 296064
rect 388438 296012 388444 296064
rect 388496 296052 388502 296064
rect 441890 296052 441896 296064
rect 388496 296024 441896 296052
rect 388496 296012 388502 296024
rect 441890 296012 441896 296024
rect 441948 296012 441954 296064
rect 372154 295944 372160 295996
rect 372212 295984 372218 295996
rect 442074 295984 442080 295996
rect 372212 295956 442080 295984
rect 372212 295944 372218 295956
rect 442074 295944 442080 295956
rect 442132 295944 442138 295996
rect 445202 295944 445208 295996
rect 445260 295984 445266 295996
rect 445260 295956 451274 295984
rect 445260 295944 445266 295956
rect 428458 295876 428464 295928
rect 428516 295916 428522 295928
rect 441706 295916 441712 295928
rect 428516 295888 441712 295916
rect 428516 295876 428522 295888
rect 441706 295876 441712 295888
rect 441764 295876 441770 295928
rect 451246 295916 451274 295956
rect 517238 295944 517244 295996
rect 517296 295984 517302 295996
rect 528830 295984 528836 295996
rect 517296 295956 528836 295984
rect 517296 295944 517302 295956
rect 528830 295944 528836 295956
rect 528888 295944 528894 295996
rect 451246 295888 513696 295916
rect 359458 295808 359464 295860
rect 359516 295848 359522 295860
rect 369854 295848 369860 295860
rect 359516 295820 369860 295848
rect 359516 295808 359522 295820
rect 369854 295808 369860 295820
rect 369912 295808 369918 295860
rect 391934 295808 391940 295860
rect 391992 295848 391998 295860
rect 393222 295848 393228 295860
rect 391992 295820 393228 295848
rect 391992 295808 391998 295820
rect 393222 295808 393228 295820
rect 393280 295848 393286 295860
rect 513558 295848 513564 295860
rect 393280 295820 513564 295848
rect 393280 295808 393286 295820
rect 513558 295808 513564 295820
rect 513616 295808 513622 295860
rect 513668 295520 513696 295888
rect 513650 295468 513656 295520
rect 513708 295468 513714 295520
rect 379238 295400 379244 295452
rect 379296 295440 379302 295452
rect 400674 295440 400680 295452
rect 379296 295412 400680 295440
rect 379296 295400 379302 295412
rect 400674 295400 400680 295412
rect 400732 295400 400738 295452
rect 302786 295332 302792 295384
rect 302844 295372 302850 295384
rect 320818 295372 320824 295384
rect 302844 295344 320824 295372
rect 302844 295332 302850 295344
rect 320818 295332 320824 295344
rect 320876 295332 320882 295384
rect 378962 295332 378968 295384
rect 379020 295372 379026 295384
rect 388438 295372 388444 295384
rect 379020 295344 388444 295372
rect 379020 295332 379026 295344
rect 388438 295332 388444 295344
rect 388496 295332 388502 295384
rect 371326 295264 371332 295316
rect 371384 295304 371390 295316
rect 378870 295304 378876 295316
rect 371384 295276 378876 295304
rect 371384 295264 371390 295276
rect 378870 295264 378876 295276
rect 378928 295264 378934 295316
rect 516134 295264 516140 295316
rect 516192 295304 516198 295316
rect 529934 295304 529940 295316
rect 516192 295276 529940 295304
rect 516192 295264 516198 295276
rect 529934 295264 529940 295276
rect 529992 295264 529998 295316
rect 371694 295196 371700 295248
rect 371752 295236 371758 295248
rect 378962 295236 378968 295248
rect 371752 295208 378968 295236
rect 371752 295196 371758 295208
rect 378962 295196 378968 295208
rect 379020 295196 379026 295248
rect 445386 295196 445392 295248
rect 445444 295236 445450 295248
rect 448606 295236 448612 295248
rect 445444 295208 448612 295236
rect 445444 295196 445450 295208
rect 448606 295196 448612 295208
rect 448664 295196 448670 295248
rect 516318 295196 516324 295248
rect 516376 295236 516382 295248
rect 528738 295236 528744 295248
rect 516376 295208 528744 295236
rect 516376 295196 516382 295208
rect 528738 295196 528744 295208
rect 528796 295196 528802 295248
rect 445478 295128 445484 295180
rect 445536 295168 445542 295180
rect 447502 295168 447508 295180
rect 445536 295140 447508 295168
rect 445536 295128 445542 295140
rect 447502 295128 447508 295140
rect 447560 295128 447566 295180
rect 516226 295128 516232 295180
rect 516284 295168 516290 295180
rect 524414 295168 524420 295180
rect 516284 295140 524420 295168
rect 516284 295128 516290 295140
rect 524414 295128 524420 295140
rect 524472 295128 524478 295180
rect 447502 294584 447508 294636
rect 447560 294624 447566 294636
rect 456058 294624 456064 294636
rect 447560 294596 456064 294624
rect 447560 294584 447566 294596
rect 456058 294584 456064 294596
rect 456116 294584 456122 294636
rect 448606 293972 448612 294024
rect 448664 294012 448670 294024
rect 449250 294012 449256 294024
rect 448664 293984 449256 294012
rect 448664 293972 448670 293984
rect 449250 293972 449256 293984
rect 449308 293972 449314 294024
rect 371234 293904 371240 293956
rect 371292 293944 371298 293956
rect 400122 293944 400128 293956
rect 371292 293916 400128 293944
rect 371292 293904 371298 293916
rect 400122 293904 400128 293916
rect 400180 293904 400186 293956
rect 516226 293904 516232 293956
rect 516284 293944 516290 293956
rect 525794 293944 525800 293956
rect 516284 293916 525800 293944
rect 516284 293904 516290 293916
rect 525794 293904 525800 293916
rect 525852 293904 525858 293956
rect 371326 293836 371332 293888
rect 371384 293876 371390 293888
rect 379238 293876 379244 293888
rect 371384 293848 379244 293876
rect 371384 293836 371390 293848
rect 379238 293836 379244 293848
rect 379296 293836 379302 293888
rect 516134 293836 516140 293888
rect 516192 293876 516198 293888
rect 523034 293876 523040 293888
rect 516192 293848 523040 293876
rect 516192 293836 516198 293848
rect 523034 293836 523040 293848
rect 523092 293836 523098 293888
rect 371234 292476 371240 292528
rect 371292 292516 371298 292528
rect 385770 292516 385776 292528
rect 371292 292488 385776 292516
rect 371292 292476 371298 292488
rect 385770 292476 385776 292488
rect 385828 292476 385834 292528
rect 516318 292476 516324 292528
rect 516376 292516 516382 292528
rect 516594 292516 516600 292528
rect 516376 292488 516600 292516
rect 516376 292476 516382 292488
rect 516594 292476 516600 292488
rect 516652 292516 516658 292528
rect 530026 292516 530032 292528
rect 516652 292488 530032 292516
rect 516652 292476 516658 292488
rect 530026 292476 530032 292488
rect 530084 292476 530090 292528
rect 516134 292408 516140 292460
rect 516192 292448 516198 292460
rect 527174 292448 527180 292460
rect 516192 292420 527180 292448
rect 516192 292408 516198 292420
rect 527174 292408 527180 292420
rect 527232 292408 527238 292460
rect 516226 292340 516232 292392
rect 516284 292380 516290 292392
rect 521654 292380 521660 292392
rect 516284 292352 521660 292380
rect 516284 292340 516290 292352
rect 521654 292340 521660 292352
rect 521712 292340 521718 292392
rect 513742 291864 513748 291916
rect 513800 291904 513806 291916
rect 514018 291904 514024 291916
rect 513800 291876 514024 291904
rect 513800 291864 513806 291876
rect 514018 291864 514024 291876
rect 514076 291864 514082 291916
rect 371694 291796 371700 291848
rect 371752 291836 371758 291848
rect 378226 291836 378232 291848
rect 371752 291808 378232 291836
rect 371752 291796 371758 291808
rect 378226 291796 378232 291808
rect 378284 291836 378290 291848
rect 379422 291836 379428 291848
rect 378284 291808 379428 291836
rect 378284 291796 378290 291808
rect 379422 291796 379428 291808
rect 379480 291796 379486 291848
rect 386322 291796 386328 291848
rect 386380 291836 386386 291848
rect 395338 291836 395344 291848
rect 386380 291808 395344 291836
rect 386380 291796 386386 291808
rect 395338 291796 395344 291808
rect 395396 291796 395402 291848
rect 372246 291728 372252 291780
rect 372304 291768 372310 291780
rect 372430 291768 372436 291780
rect 372304 291740 372436 291768
rect 372304 291728 372310 291740
rect 372430 291728 372436 291740
rect 372488 291728 372494 291780
rect 371694 291184 371700 291236
rect 371752 291224 371758 291236
rect 385678 291224 385684 291236
rect 371752 291196 385684 291224
rect 371752 291184 371758 291196
rect 385678 291184 385684 291196
rect 385736 291224 385742 291236
rect 386322 291224 386328 291236
rect 385736 291196 386328 291224
rect 385736 291184 385742 291196
rect 386322 291184 386328 291196
rect 386380 291184 386386 291236
rect 380894 291116 380900 291168
rect 380952 291156 380958 291168
rect 382182 291156 382188 291168
rect 380952 291128 382188 291156
rect 380952 291116 380958 291128
rect 382182 291116 382188 291128
rect 382240 291116 382246 291168
rect 516318 291116 516324 291168
rect 516376 291156 516382 291168
rect 516778 291156 516784 291168
rect 516376 291128 516784 291156
rect 516376 291116 516382 291128
rect 516778 291116 516784 291128
rect 516836 291156 516842 291168
rect 530118 291156 530124 291168
rect 516836 291128 530124 291156
rect 516836 291116 516842 291128
rect 530118 291116 530124 291128
rect 530176 291116 530182 291168
rect 516226 291048 516232 291100
rect 516284 291088 516290 291100
rect 516686 291088 516692 291100
rect 516284 291060 516692 291088
rect 516284 291048 516290 291060
rect 516686 291048 516692 291060
rect 516744 291088 516750 291100
rect 528646 291088 528652 291100
rect 516744 291060 528652 291088
rect 516744 291048 516750 291060
rect 528646 291048 528652 291060
rect 528704 291048 528710 291100
rect 371326 290640 371332 290692
rect 371384 290680 371390 290692
rect 371878 290680 371884 290692
rect 371384 290652 371884 290680
rect 371384 290640 371390 290652
rect 371878 290640 371884 290652
rect 371936 290640 371942 290692
rect 371694 290504 371700 290556
rect 371752 290544 371758 290556
rect 380894 290544 380900 290556
rect 371752 290516 380900 290544
rect 371752 290504 371758 290516
rect 380894 290504 380900 290516
rect 380952 290504 380958 290556
rect 371786 290436 371792 290488
rect 371844 290476 371850 290488
rect 382274 290476 382280 290488
rect 371844 290448 382280 290476
rect 371844 290436 371850 290448
rect 382274 290436 382280 290448
rect 382332 290436 382338 290488
rect 445478 290368 445484 290420
rect 445536 290408 445542 290420
rect 447410 290408 447416 290420
rect 445536 290380 447416 290408
rect 445536 290368 445542 290380
rect 447410 290368 447416 290380
rect 447468 290408 447474 290420
rect 447962 290408 447968 290420
rect 447468 290380 447968 290408
rect 447468 290368 447474 290380
rect 447962 290368 447968 290380
rect 448020 290368 448026 290420
rect 170398 289824 170404 289876
rect 170456 289864 170462 289876
rect 197354 289864 197360 289876
rect 170456 289836 197360 289864
rect 170456 289824 170462 289836
rect 197354 289824 197360 289836
rect 197412 289824 197418 289876
rect 444282 289824 444288 289876
rect 444340 289864 444346 289876
rect 447870 289864 447876 289876
rect 444340 289836 447876 289864
rect 444340 289824 444346 289836
rect 447870 289824 447876 289836
rect 447928 289824 447934 289876
rect 376018 289756 376024 289808
rect 376076 289796 376082 289808
rect 377398 289796 377404 289808
rect 376076 289768 377404 289796
rect 376076 289756 376082 289768
rect 377398 289756 377404 289768
rect 377456 289756 377462 289808
rect 378134 289756 378140 289808
rect 378192 289796 378198 289808
rect 378778 289796 378784 289808
rect 378192 289768 378784 289796
rect 378192 289756 378198 289768
rect 378778 289756 378784 289768
rect 378836 289756 378842 289808
rect 516318 289756 516324 289808
rect 516376 289796 516382 289808
rect 516502 289796 516508 289808
rect 516376 289768 516508 289796
rect 516376 289756 516382 289768
rect 516502 289756 516508 289768
rect 516560 289796 516566 289808
rect 528554 289796 528560 289808
rect 516560 289768 528560 289796
rect 516560 289756 516566 289768
rect 528554 289756 528560 289768
rect 528612 289756 528618 289808
rect 516226 289688 516232 289740
rect 516284 289728 516290 289740
rect 525886 289728 525892 289740
rect 516284 289700 525892 289728
rect 516284 289688 516290 289700
rect 525886 289688 525892 289700
rect 525944 289688 525950 289740
rect 516134 289620 516140 289672
rect 516192 289660 516198 289672
rect 524506 289660 524512 289672
rect 516192 289632 524512 289660
rect 516192 289620 516198 289632
rect 524506 289620 524512 289632
rect 524564 289620 524570 289672
rect 302234 289212 302240 289264
rect 302292 289252 302298 289264
rect 304350 289252 304356 289264
rect 302292 289224 304356 289252
rect 302292 289212 302298 289224
rect 304350 289212 304356 289224
rect 304408 289212 304414 289264
rect 371694 289212 371700 289264
rect 371752 289252 371758 289264
rect 376018 289252 376024 289264
rect 371752 289224 376024 289252
rect 371752 289212 371758 289224
rect 376018 289212 376024 289224
rect 376076 289212 376082 289264
rect 371234 289076 371240 289128
rect 371292 289116 371298 289128
rect 378134 289116 378140 289128
rect 371292 289088 378140 289116
rect 371292 289076 371298 289088
rect 378134 289076 378140 289088
rect 378192 289076 378198 289128
rect 371694 288532 371700 288584
rect 371752 288572 371758 288584
rect 375926 288572 375932 288584
rect 371752 288544 375932 288572
rect 371752 288532 371758 288544
rect 375926 288532 375932 288544
rect 375984 288532 375990 288584
rect 445938 287444 445944 287496
rect 445996 287484 446002 287496
rect 446674 287484 446680 287496
rect 445996 287456 446680 287484
rect 445996 287444 446002 287456
rect 446674 287444 446680 287456
rect 446732 287444 446738 287496
rect 443178 287104 443184 287156
rect 443236 287144 443242 287156
rect 447778 287144 447784 287156
rect 443236 287116 447784 287144
rect 443236 287104 443242 287116
rect 447778 287104 447784 287116
rect 447836 287104 447842 287156
rect 178678 287036 178684 287088
rect 178736 287076 178742 287088
rect 198550 287076 198556 287088
rect 178736 287048 198556 287076
rect 178736 287036 178742 287048
rect 198550 287036 198556 287048
rect 198608 287036 198614 287088
rect 302234 286492 302240 286544
rect 302292 286532 302298 286544
rect 304258 286532 304264 286544
rect 302292 286504 304264 286532
rect 302292 286492 302298 286504
rect 304258 286492 304264 286504
rect 304316 286492 304322 286544
rect 371142 286356 371148 286408
rect 371200 286396 371206 286408
rect 371602 286396 371608 286408
rect 371200 286368 371608 286396
rect 371200 286356 371206 286368
rect 371602 286356 371608 286368
rect 371660 286356 371666 286408
rect 371510 286288 371516 286340
rect 371568 286328 371574 286340
rect 377398 286328 377404 286340
rect 371568 286300 377404 286328
rect 371568 286288 371574 286300
rect 377398 286288 377404 286300
rect 377456 286288 377462 286340
rect 371970 285676 371976 285728
rect 372028 285716 372034 285728
rect 374546 285716 374552 285728
rect 372028 285688 374552 285716
rect 372028 285676 372034 285688
rect 374546 285676 374552 285688
rect 374604 285676 374610 285728
rect 444742 284792 444748 284844
rect 444800 284832 444806 284844
rect 446398 284832 446404 284844
rect 444800 284804 446404 284832
rect 444800 284792 444806 284804
rect 446398 284792 446404 284804
rect 446456 284792 446462 284844
rect 372246 284316 372252 284368
rect 372304 284356 372310 284368
rect 375374 284356 375380 284368
rect 372304 284328 375380 284356
rect 372304 284316 372310 284328
rect 375374 284316 375380 284328
rect 375432 284316 375438 284368
rect 369210 283568 369216 283620
rect 369268 283608 369274 283620
rect 369670 283608 369676 283620
rect 369268 283580 369676 283608
rect 369268 283568 369274 283580
rect 369670 283568 369676 283580
rect 369728 283568 369734 283620
rect 371510 283568 371516 283620
rect 371568 283608 371574 283620
rect 376754 283608 376760 283620
rect 371568 283580 376760 283608
rect 371568 283568 371574 283580
rect 376754 283568 376760 283580
rect 376812 283608 376818 283620
rect 376938 283608 376944 283620
rect 376812 283580 376944 283608
rect 376812 283568 376818 283580
rect 376938 283568 376944 283580
rect 376996 283568 377002 283620
rect 369118 283296 369124 283348
rect 369176 283336 369182 283348
rect 369394 283336 369400 283348
rect 369176 283308 369400 283336
rect 369176 283296 369182 283308
rect 369394 283296 369400 283308
rect 369452 283296 369458 283348
rect 174538 282888 174544 282940
rect 174596 282928 174602 282940
rect 197354 282928 197360 282940
rect 174596 282900 197360 282928
rect 174596 282888 174602 282900
rect 197354 282888 197360 282900
rect 197412 282888 197418 282940
rect 302786 282888 302792 282940
rect 302844 282928 302850 282940
rect 353938 282928 353944 282940
rect 302844 282900 353944 282928
rect 302844 282888 302850 282900
rect 353938 282888 353944 282900
rect 353996 282888 354002 282940
rect 445846 282888 445852 282940
rect 445904 282928 445910 282940
rect 446582 282928 446588 282940
rect 445904 282900 446588 282928
rect 445904 282888 445910 282900
rect 446582 282888 446588 282900
rect 446640 282888 446646 282940
rect 377582 282820 377588 282872
rect 377640 282860 377646 282872
rect 378042 282860 378048 282872
rect 377640 282832 378048 282860
rect 377640 282820 377646 282832
rect 378042 282820 378048 282832
rect 378100 282860 378106 282872
rect 425698 282860 425704 282872
rect 378100 282832 425704 282860
rect 378100 282820 378106 282832
rect 425698 282820 425704 282832
rect 425756 282820 425762 282872
rect 444374 282820 444380 282872
rect 444432 282860 444438 282872
rect 446214 282860 446220 282872
rect 444432 282832 446220 282860
rect 444432 282820 444438 282832
rect 446214 282820 446220 282832
rect 446272 282820 446278 282872
rect 371694 282276 371700 282328
rect 371752 282316 371758 282328
rect 375466 282316 375472 282328
rect 371752 282288 375472 282316
rect 371752 282276 371758 282288
rect 375466 282276 375472 282288
rect 375524 282316 375530 282328
rect 377674 282316 377680 282328
rect 375524 282288 377680 282316
rect 375524 282276 375530 282288
rect 377674 282276 377680 282288
rect 377732 282276 377738 282328
rect 371602 282208 371608 282260
rect 371660 282248 371666 282260
rect 375834 282248 375840 282260
rect 371660 282220 375840 282248
rect 371660 282208 371666 282220
rect 375834 282208 375840 282220
rect 375892 282248 375898 282260
rect 376846 282248 376852 282260
rect 375892 282220 376852 282248
rect 375892 282208 375898 282220
rect 376846 282208 376852 282220
rect 376904 282208 376910 282260
rect 371510 282140 371516 282192
rect 371568 282180 371574 282192
rect 378042 282180 378048 282192
rect 371568 282152 378048 282180
rect 371568 282140 371574 282152
rect 378042 282140 378048 282152
rect 378100 282140 378106 282192
rect 160094 281528 160100 281580
rect 160152 281568 160158 281580
rect 197906 281568 197912 281580
rect 160152 281540 197912 281568
rect 160152 281528 160158 281540
rect 197906 281528 197912 281540
rect 197964 281528 197970 281580
rect 516134 281528 516140 281580
rect 516192 281568 516198 281580
rect 524506 281568 524512 281580
rect 516192 281540 524512 281568
rect 516192 281528 516198 281540
rect 524506 281528 524512 281540
rect 524564 281528 524570 281580
rect 377490 281460 377496 281512
rect 377548 281500 377554 281512
rect 378042 281500 378048 281512
rect 377548 281472 378048 281500
rect 377548 281460 377554 281472
rect 378042 281460 378048 281472
rect 378100 281500 378106 281512
rect 428458 281500 428464 281512
rect 378100 281472 428464 281500
rect 378100 281460 378106 281472
rect 428458 281460 428464 281472
rect 428516 281460 428522 281512
rect 444742 281256 444748 281308
rect 444800 281296 444806 281308
rect 445754 281296 445760 281308
rect 444800 281268 445760 281296
rect 444800 281256 444806 281268
rect 445754 281256 445760 281268
rect 445812 281296 445818 281308
rect 446766 281296 446772 281308
rect 445812 281268 446772 281296
rect 445812 281256 445818 281268
rect 446766 281256 446772 281268
rect 446824 281256 446830 281308
rect 369210 280848 369216 280900
rect 369268 280888 369274 280900
rect 369394 280888 369400 280900
rect 369268 280860 369400 280888
rect 369268 280848 369274 280860
rect 369394 280848 369400 280860
rect 369452 280848 369458 280900
rect 371510 280780 371516 280832
rect 371568 280820 371574 280832
rect 378042 280820 378048 280832
rect 371568 280792 378048 280820
rect 371568 280780 371574 280792
rect 378042 280780 378048 280792
rect 378100 280780 378106 280832
rect 445478 280576 445484 280628
rect 445536 280616 445542 280628
rect 447318 280616 447324 280628
rect 445536 280588 447324 280616
rect 445536 280576 445542 280588
rect 447318 280576 447324 280588
rect 447376 280616 447382 280628
rect 448054 280616 448060 280628
rect 447376 280588 448060 280616
rect 447376 280576 447382 280588
rect 448054 280576 448060 280588
rect 448112 280576 448118 280628
rect 516134 280440 516140 280492
rect 516192 280480 516198 280492
rect 518894 280480 518900 280492
rect 516192 280452 518900 280480
rect 516192 280440 516198 280452
rect 518894 280440 518900 280452
rect 518952 280440 518958 280492
rect 516226 280168 516232 280220
rect 516284 280208 516290 280220
rect 521654 280208 521660 280220
rect 516284 280180 521660 280208
rect 516284 280168 516290 280180
rect 521654 280168 521660 280180
rect 521712 280168 521718 280220
rect 371418 279420 371424 279472
rect 371476 279460 371482 279472
rect 377030 279460 377036 279472
rect 371476 279432 377036 279460
rect 371476 279420 371482 279432
rect 377030 279420 377036 279432
rect 377088 279420 377094 279472
rect 517790 279420 517796 279472
rect 517848 279460 517854 279472
rect 521930 279460 521936 279472
rect 517848 279432 521936 279460
rect 517848 279420 517854 279432
rect 521930 279420 521936 279432
rect 521988 279420 521994 279472
rect 371602 279352 371608 279404
rect 371660 279392 371666 279404
rect 373994 279392 374000 279404
rect 371660 279364 374000 279392
rect 371660 279352 371666 279364
rect 373994 279352 374000 279364
rect 374052 279392 374058 279404
rect 374730 279392 374736 279404
rect 374052 279364 374736 279392
rect 374052 279352 374058 279364
rect 374730 279352 374736 279364
rect 374788 279352 374794 279404
rect 516134 278808 516140 278860
rect 516192 278848 516198 278860
rect 523126 278848 523132 278860
rect 516192 278820 523132 278848
rect 516192 278808 516198 278820
rect 523126 278808 523132 278820
rect 523184 278808 523190 278860
rect 175918 278740 175924 278792
rect 175976 278780 175982 278792
rect 197538 278780 197544 278792
rect 175976 278752 197544 278780
rect 175976 278740 175982 278752
rect 197538 278740 197544 278752
rect 197596 278740 197602 278792
rect 302418 278740 302424 278792
rect 302476 278780 302482 278792
rect 356698 278780 356704 278792
rect 302476 278752 356704 278780
rect 302476 278740 302482 278752
rect 356698 278740 356704 278752
rect 356756 278740 356762 278792
rect 516226 278740 516232 278792
rect 516284 278780 516290 278792
rect 524414 278780 524420 278792
rect 516284 278752 524420 278780
rect 516284 278740 516290 278752
rect 524414 278740 524420 278752
rect 524472 278740 524478 278792
rect 376110 278672 376116 278724
rect 376168 278712 376174 278724
rect 377030 278712 377036 278724
rect 376168 278684 377036 278712
rect 376168 278672 376174 278684
rect 377030 278672 377036 278684
rect 377088 278672 377094 278724
rect 516134 278672 516140 278724
rect 516192 278712 516198 278724
rect 516410 278712 516416 278724
rect 516192 278684 516416 278712
rect 516192 278672 516198 278684
rect 516410 278672 516416 278684
rect 516468 278672 516474 278724
rect 371602 278264 371608 278316
rect 371660 278304 371666 278316
rect 374086 278304 374092 278316
rect 371660 278276 374092 278304
rect 371660 278264 371666 278276
rect 374086 278264 374092 278276
rect 374144 278304 374150 278316
rect 374822 278304 374828 278316
rect 374144 278276 374828 278304
rect 374144 278264 374150 278276
rect 374822 278264 374828 278276
rect 374880 278264 374886 278316
rect 516686 277856 516692 277908
rect 516744 277896 516750 277908
rect 518250 277896 518256 277908
rect 516744 277868 518256 277896
rect 516744 277856 516750 277868
rect 518250 277856 518256 277868
rect 518308 277856 518314 277908
rect 518250 277448 518256 277500
rect 518308 277488 518314 277500
rect 519262 277488 519268 277500
rect 518308 277460 519268 277488
rect 518308 277448 518314 277460
rect 519262 277448 519268 277460
rect 519320 277448 519326 277500
rect 181438 277380 181444 277432
rect 181496 277420 181502 277432
rect 197354 277420 197360 277432
rect 181496 277392 197360 277420
rect 181496 277380 181502 277392
rect 197354 277380 197360 277392
rect 197412 277380 197418 277432
rect 516410 277380 516416 277432
rect 516468 277420 516474 277432
rect 521746 277420 521752 277432
rect 516468 277392 521752 277420
rect 516468 277380 516474 277392
rect 521746 277380 521752 277392
rect 521804 277380 521810 277432
rect 516134 276904 516140 276956
rect 516192 276944 516198 276956
rect 516410 276944 516416 276956
rect 516192 276916 516416 276944
rect 516192 276904 516198 276916
rect 516410 276904 516416 276916
rect 516468 276904 516474 276956
rect 516134 276768 516140 276820
rect 516192 276808 516198 276820
rect 519170 276808 519176 276820
rect 516192 276780 519176 276808
rect 516192 276768 516198 276780
rect 519170 276768 519176 276780
rect 519228 276768 519234 276820
rect 516686 276292 516692 276344
rect 516744 276332 516750 276344
rect 518066 276332 518072 276344
rect 516744 276304 518072 276332
rect 516744 276292 516750 276304
rect 518066 276292 518072 276304
rect 518124 276332 518130 276344
rect 520274 276332 520280 276344
rect 518124 276304 520280 276332
rect 518124 276292 518130 276304
rect 520274 276292 520280 276304
rect 520332 276292 520338 276344
rect 372430 276224 372436 276276
rect 372488 276264 372494 276276
rect 373902 276264 373908 276276
rect 372488 276236 373908 276264
rect 372488 276224 372494 276236
rect 373902 276224 373908 276236
rect 373960 276224 373966 276276
rect 371418 276156 371424 276208
rect 371476 276196 371482 276208
rect 374638 276196 374644 276208
rect 371476 276168 374644 276196
rect 371476 276156 371482 276168
rect 374638 276156 374644 276168
rect 374696 276156 374702 276208
rect 519170 276088 519176 276140
rect 519228 276128 519234 276140
rect 520458 276128 520464 276140
rect 519228 276100 520464 276128
rect 519228 276088 519234 276100
rect 520458 276088 520464 276100
rect 520516 276088 520522 276140
rect 302786 276020 302792 276072
rect 302844 276060 302850 276072
rect 358170 276060 358176 276072
rect 302844 276032 358176 276060
rect 302844 276020 302850 276032
rect 358170 276020 358176 276032
rect 358228 276020 358234 276072
rect 516318 276020 516324 276072
rect 516376 276060 516382 276072
rect 521930 276060 521936 276072
rect 516376 276032 521936 276060
rect 516376 276020 516382 276032
rect 521930 276020 521936 276032
rect 521988 276020 521994 276072
rect 371602 275748 371608 275800
rect 371660 275788 371666 275800
rect 374178 275788 374184 275800
rect 371660 275760 374184 275788
rect 371660 275748 371666 275760
rect 374178 275748 374184 275760
rect 374236 275748 374242 275800
rect 372798 275340 372804 275392
rect 372856 275380 372862 275392
rect 373258 275380 373264 275392
rect 372856 275352 373264 275380
rect 372856 275340 372862 275352
rect 373258 275340 373264 275352
rect 373316 275340 373322 275392
rect 372154 275204 372160 275256
rect 372212 275244 372218 275256
rect 373258 275244 373264 275256
rect 372212 275216 373264 275244
rect 372212 275204 372218 275216
rect 373258 275204 373264 275216
rect 373316 275244 373322 275256
rect 374270 275244 374276 275256
rect 373316 275216 374276 275244
rect 373316 275204 373322 275216
rect 374270 275204 374276 275216
rect 374328 275204 374334 275256
rect 516134 275204 516140 275256
rect 516192 275244 516198 275256
rect 519078 275244 519084 275256
rect 516192 275216 519084 275244
rect 516192 275204 516198 275216
rect 519078 275204 519084 275216
rect 519136 275204 519142 275256
rect 516318 275136 516324 275188
rect 516376 275176 516382 275188
rect 520550 275176 520556 275188
rect 516376 275148 520556 275176
rect 516376 275136 516382 275148
rect 520550 275136 520556 275148
rect 520608 275136 520614 275188
rect 188338 274660 188344 274712
rect 188396 274700 188402 274712
rect 197538 274700 197544 274712
rect 188396 274672 197544 274700
rect 188396 274660 188402 274672
rect 197538 274660 197544 274672
rect 197596 274660 197602 274712
rect 516134 274660 516140 274712
rect 516192 274700 516198 274712
rect 518342 274700 518348 274712
rect 516192 274672 518348 274700
rect 516192 274660 516198 274672
rect 518342 274660 518348 274672
rect 518400 274660 518406 274712
rect 373350 274592 373356 274644
rect 373408 274632 373414 274644
rect 374178 274632 374184 274644
rect 373408 274604 374184 274632
rect 373408 274592 373414 274604
rect 374178 274592 374184 274604
rect 374236 274592 374242 274644
rect 516686 274048 516692 274100
rect 516744 274088 516750 274100
rect 517606 274088 517612 274100
rect 516744 274060 517612 274088
rect 516744 274048 516750 274060
rect 517606 274048 517612 274060
rect 517664 274088 517670 274100
rect 519170 274088 519176 274100
rect 517664 274060 519176 274088
rect 517664 274048 517670 274060
rect 519170 274048 519176 274060
rect 519228 274048 519234 274100
rect 371602 273572 371608 273624
rect 371660 273612 371666 273624
rect 373994 273612 374000 273624
rect 371660 273584 374000 273612
rect 371660 273572 371666 273584
rect 373994 273572 374000 273584
rect 374052 273612 374058 273624
rect 374362 273612 374368 273624
rect 374052 273584 374368 273612
rect 374052 273572 374058 273584
rect 374362 273572 374368 273584
rect 374420 273572 374426 273624
rect 180058 273232 180064 273284
rect 180116 273272 180122 273284
rect 197354 273272 197360 273284
rect 180116 273244 197360 273272
rect 180116 273232 180122 273244
rect 197354 273232 197360 273244
rect 197412 273232 197418 273284
rect 302694 273232 302700 273284
rect 302752 273272 302758 273284
rect 360562 273272 360568 273284
rect 302752 273244 360568 273272
rect 302752 273232 302758 273244
rect 360562 273232 360568 273244
rect 360620 273232 360626 273284
rect 371510 273232 371516 273284
rect 371568 273272 371574 273284
rect 372614 273272 372620 273284
rect 371568 273244 372620 273272
rect 371568 273232 371574 273244
rect 372614 273232 372620 273244
rect 372672 273272 372678 273284
rect 372890 273272 372896 273284
rect 372672 273244 372896 273272
rect 372672 273232 372678 273244
rect 372890 273232 372896 273244
rect 372948 273232 372954 273284
rect 517514 273232 517520 273284
rect 517572 273272 517578 273284
rect 518250 273272 518256 273284
rect 517572 273244 518256 273272
rect 517572 273232 517578 273244
rect 518250 273232 518256 273244
rect 518308 273232 518314 273284
rect 444558 273164 444564 273216
rect 444616 273204 444622 273216
rect 447134 273204 447140 273216
rect 444616 273176 447140 273204
rect 444616 273164 444622 273176
rect 447134 273164 447140 273176
rect 447192 273164 447198 273216
rect 516134 273164 516140 273216
rect 516192 273204 516198 273216
rect 524782 273204 524788 273216
rect 516192 273176 524788 273204
rect 516192 273164 516198 273176
rect 524782 273164 524788 273176
rect 524840 273204 524846 273216
rect 528646 273204 528652 273216
rect 524840 273176 528652 273204
rect 524840 273164 524846 273176
rect 528646 273164 528652 273176
rect 528704 273164 528710 273216
rect 516318 272484 516324 272536
rect 516376 272524 516382 272536
rect 517882 272524 517888 272536
rect 516376 272496 517888 272524
rect 516376 272484 516382 272496
rect 517882 272484 517888 272496
rect 517940 272484 517946 272536
rect 516134 271872 516140 271924
rect 516192 271912 516198 271924
rect 525886 271912 525892 271924
rect 516192 271884 525892 271912
rect 516192 271872 516198 271884
rect 525886 271872 525892 271884
rect 525944 271872 525950 271924
rect 371878 271804 371884 271856
rect 371936 271844 371942 271856
rect 372246 271844 372252 271856
rect 371936 271816 372252 271844
rect 371936 271804 371942 271816
rect 372246 271804 372252 271816
rect 372304 271844 372310 271856
rect 377214 271844 377220 271856
rect 372304 271816 377220 271844
rect 372304 271804 372310 271816
rect 377214 271804 377220 271816
rect 377272 271804 377278 271856
rect 371694 271736 371700 271788
rect 371752 271776 371758 271788
rect 377122 271776 377128 271788
rect 371752 271748 377128 271776
rect 371752 271736 371758 271748
rect 377122 271736 377128 271748
rect 377180 271736 377186 271788
rect 371786 271668 371792 271720
rect 371844 271708 371850 271720
rect 372154 271708 372160 271720
rect 371844 271680 372160 271708
rect 371844 271668 371850 271680
rect 372154 271668 372160 271680
rect 372212 271708 372218 271720
rect 376202 271708 376208 271720
rect 372212 271680 376208 271708
rect 372212 271668 372218 271680
rect 376202 271668 376208 271680
rect 376260 271668 376266 271720
rect 516134 271192 516140 271244
rect 516192 271232 516198 271244
rect 521010 271232 521016 271244
rect 516192 271204 521016 271232
rect 516192 271192 516198 271204
rect 521010 271192 521016 271204
rect 521068 271232 521074 271244
rect 524598 271232 524604 271244
rect 521068 271204 524604 271232
rect 521068 271192 521074 271204
rect 524598 271192 524604 271204
rect 524656 271192 524662 271244
rect 516318 271124 516324 271176
rect 516376 271164 516382 271176
rect 521838 271164 521844 271176
rect 516376 271136 521844 271164
rect 516376 271124 516382 271136
rect 521838 271124 521844 271136
rect 521896 271164 521902 271176
rect 522022 271164 522028 271176
rect 521896 271136 522028 271164
rect 521896 271124 521902 271136
rect 522022 271124 522028 271136
rect 522080 271124 522086 271176
rect 372522 270580 372528 270632
rect 372580 270620 372586 270632
rect 375558 270620 375564 270632
rect 372580 270592 375564 270620
rect 372580 270580 372586 270592
rect 375558 270580 375564 270592
rect 375616 270580 375622 270632
rect 186958 270512 186964 270564
rect 187016 270552 187022 270564
rect 197538 270552 197544 270564
rect 187016 270524 197544 270552
rect 187016 270512 187022 270524
rect 197538 270512 197544 270524
rect 197596 270512 197602 270564
rect 371786 270444 371792 270496
rect 371844 270484 371850 270496
rect 372062 270484 372068 270496
rect 371844 270456 372068 270484
rect 371844 270444 371850 270456
rect 372062 270444 372068 270456
rect 372120 270484 372126 270496
rect 374454 270484 374460 270496
rect 372120 270456 374460 270484
rect 372120 270444 372126 270456
rect 374454 270444 374460 270456
rect 374512 270444 374518 270496
rect 516134 270172 516140 270224
rect 516192 270212 516198 270224
rect 519630 270212 519636 270224
rect 516192 270184 519636 270212
rect 516192 270172 516198 270184
rect 519630 270172 519636 270184
rect 519688 270212 519694 270224
rect 523034 270212 523040 270224
rect 519688 270184 523040 270212
rect 519688 270172 519694 270184
rect 523034 270172 523040 270184
rect 523092 270172 523098 270224
rect 377306 270076 377312 270088
rect 373966 270048 377312 270076
rect 371418 269764 371424 269816
rect 371476 269804 371482 269816
rect 373966 269804 373994 270048
rect 377306 270036 377312 270048
rect 377364 270076 377370 270088
rect 441614 270076 441620 270088
rect 377364 270048 441620 270076
rect 377364 270036 377370 270048
rect 441614 270036 441620 270048
rect 441672 270036 441678 270088
rect 371476 269776 373994 269804
rect 371476 269764 371482 269776
rect 445478 269764 445484 269816
rect 445536 269804 445542 269816
rect 447226 269804 447232 269816
rect 445536 269776 447232 269804
rect 445536 269764 445542 269776
rect 447226 269764 447232 269776
rect 447284 269764 447290 269816
rect 516318 269492 516324 269544
rect 516376 269532 516382 269544
rect 520642 269532 520648 269544
rect 516376 269504 520648 269532
rect 516376 269492 516382 269504
rect 520642 269492 520648 269504
rect 520700 269492 520706 269544
rect 193858 269288 193864 269340
rect 193916 269328 193922 269340
rect 198458 269328 198464 269340
rect 193916 269300 198464 269328
rect 193916 269288 193922 269300
rect 198458 269288 198464 269300
rect 198516 269288 198522 269340
rect 516134 269084 516140 269136
rect 516192 269124 516198 269136
rect 525794 269124 525800 269136
rect 516192 269096 525800 269124
rect 516192 269084 516198 269096
rect 525794 269084 525800 269096
rect 525852 269084 525858 269136
rect 371878 269016 371884 269068
rect 371936 269056 371942 269068
rect 375650 269056 375656 269068
rect 371936 269028 375656 269056
rect 371936 269016 371942 269028
rect 375650 269016 375656 269028
rect 375708 269016 375714 269068
rect 471054 269016 471060 269068
rect 471112 269056 471118 269068
rect 471238 269056 471244 269068
rect 471112 269028 471244 269056
rect 471112 269016 471118 269028
rect 471238 269016 471244 269028
rect 471296 269056 471302 269068
rect 513374 269056 513380 269068
rect 471296 269028 513380 269056
rect 471296 269016 471302 269028
rect 513374 269016 513380 269028
rect 513432 269016 513438 269068
rect 371970 268948 371976 269000
rect 372028 268988 372034 269000
rect 373074 268988 373080 269000
rect 372028 268960 373080 268988
rect 372028 268948 372034 268960
rect 373074 268948 373080 268960
rect 373132 268948 373138 269000
rect 513282 268948 513288 269000
rect 513340 268988 513346 269000
rect 514754 268988 514760 269000
rect 513340 268960 514760 268988
rect 513340 268948 513346 268960
rect 514754 268948 514760 268960
rect 514812 268948 514818 269000
rect 516134 268608 516140 268660
rect 516192 268648 516198 268660
rect 520366 268648 520372 268660
rect 516192 268620 520372 268648
rect 516192 268608 516198 268620
rect 520366 268608 520372 268620
rect 520424 268608 520430 268660
rect 486418 268540 486424 268592
rect 486476 268580 486482 268592
rect 516502 268580 516508 268592
rect 486476 268552 516508 268580
rect 486476 268540 486482 268552
rect 516502 268540 516508 268552
rect 516560 268540 516566 268592
rect 445478 268472 445484 268524
rect 445536 268512 445542 268524
rect 445754 268512 445760 268524
rect 445536 268484 445760 268512
rect 445536 268472 445542 268484
rect 445754 268472 445760 268484
rect 445812 268512 445818 268524
rect 471054 268512 471060 268524
rect 445812 268484 471060 268512
rect 445812 268472 445818 268484
rect 471054 268472 471060 268484
rect 471112 268472 471118 268524
rect 476758 268472 476764 268524
rect 476816 268512 476822 268524
rect 516410 268512 516416 268524
rect 476816 268484 516416 268512
rect 476816 268472 476822 268484
rect 516410 268472 516416 268484
rect 516468 268472 516474 268524
rect 303338 268404 303344 268456
rect 303396 268444 303402 268456
rect 369946 268444 369952 268456
rect 303396 268416 369952 268444
rect 303396 268404 303402 268416
rect 369946 268404 369952 268416
rect 370004 268404 370010 268456
rect 457438 268404 457444 268456
rect 457496 268444 457502 268456
rect 516594 268444 516600 268456
rect 457496 268416 516600 268444
rect 457496 268404 457502 268416
rect 516594 268404 516600 268416
rect 516652 268404 516658 268456
rect 303246 268336 303252 268388
rect 303304 268376 303310 268388
rect 370682 268376 370688 268388
rect 303304 268348 370688 268376
rect 303304 268336 303310 268348
rect 370682 268336 370688 268348
rect 370740 268336 370746 268388
rect 444558 268336 444564 268388
rect 444616 268376 444622 268388
rect 445478 268376 445484 268388
rect 444616 268348 445484 268376
rect 444616 268336 444622 268348
rect 445478 268336 445484 268348
rect 445536 268336 445542 268388
rect 449342 268336 449348 268388
rect 449400 268376 449406 268388
rect 516778 268376 516784 268388
rect 449400 268348 516784 268376
rect 449400 268336 449406 268348
rect 516778 268336 516784 268348
rect 516836 268336 516842 268388
rect 369946 268268 369952 268320
rect 370004 268308 370010 268320
rect 370222 268308 370228 268320
rect 370004 268280 370228 268308
rect 370004 268268 370010 268280
rect 370222 268268 370228 268280
rect 370280 268268 370286 268320
rect 369118 268200 369124 268252
rect 369176 268200 369182 268252
rect 369026 267996 369032 268048
rect 369084 268036 369090 268048
rect 369136 268036 369164 268200
rect 369084 268008 369164 268036
rect 369084 267996 369090 268008
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 10318 267696 10324 267708
rect 3016 267668 10324 267696
rect 3016 267656 3022 267668
rect 10318 267656 10324 267668
rect 10376 267656 10382 267708
rect 449158 267656 449164 267708
rect 449216 267696 449222 267708
rect 516226 267696 516232 267708
rect 449216 267668 516232 267696
rect 449216 267656 449222 267668
rect 516226 267656 516232 267668
rect 516284 267656 516290 267708
rect 303154 266976 303160 267028
rect 303212 267016 303218 267028
rect 370590 267016 370596 267028
rect 303212 266988 370596 267016
rect 303212 266976 303218 266988
rect 370590 266976 370596 266988
rect 370648 266976 370654 267028
rect 184198 266364 184204 266416
rect 184256 266404 184262 266416
rect 197630 266404 197636 266416
rect 184256 266376 197636 266404
rect 184256 266364 184262 266376
rect 197630 266364 197636 266376
rect 197688 266364 197694 266416
rect 362862 266296 362868 266348
rect 362920 266336 362926 266348
rect 431770 266336 431776 266348
rect 362920 266308 431776 266336
rect 362920 266296 362926 266308
rect 431770 266296 431776 266308
rect 431828 266336 431834 266348
rect 434898 266336 434904 266348
rect 431828 266308 434904 266336
rect 431828 266296 431834 266308
rect 434898 266296 434904 266308
rect 434956 266336 434962 266348
rect 434956 266308 503668 266336
rect 434956 266296 434962 266308
rect 364886 266228 364892 266280
rect 364944 266268 364950 266280
rect 431862 266268 431868 266280
rect 364944 266240 431868 266268
rect 364944 266228 364950 266240
rect 431862 266228 431868 266240
rect 431920 266268 431926 266280
rect 436922 266268 436928 266280
rect 431920 266240 436928 266268
rect 431920 266228 431926 266240
rect 436922 266228 436928 266240
rect 436980 266268 436986 266280
rect 503640 266268 503668 266308
rect 503714 266296 503720 266348
rect 503772 266336 503778 266348
rect 504910 266336 504916 266348
rect 503772 266308 504916 266336
rect 503772 266296 503778 266308
rect 504910 266296 504916 266308
rect 504968 266296 504974 266348
rect 506842 266296 506848 266348
rect 506900 266336 506906 266348
rect 507762 266336 507768 266348
rect 506900 266308 507768 266336
rect 506900 266296 506906 266308
rect 507762 266296 507768 266308
rect 507820 266336 507826 266348
rect 513742 266336 513748 266348
rect 507820 266308 513748 266336
rect 507820 266296 507826 266308
rect 513742 266296 513748 266308
rect 513800 266296 513806 266348
rect 506860 266268 506888 266296
rect 436980 266240 489914 266268
rect 503640 266240 506888 266268
rect 436980 266228 436986 266240
rect 353938 266160 353944 266212
rect 353996 266200 354002 266212
rect 368934 266200 368940 266212
rect 353996 266172 368940 266200
rect 353996 266160 354002 266172
rect 368934 266160 368940 266172
rect 368992 266200 368998 266212
rect 369118 266200 369124 266212
rect 368992 266172 369124 266200
rect 368992 266160 368998 266172
rect 369118 266160 369124 266172
rect 369176 266200 369182 266212
rect 370222 266200 370228 266212
rect 369176 266172 370228 266200
rect 369176 266160 369182 266172
rect 370222 266160 370228 266172
rect 370280 266160 370286 266212
rect 429838 266160 429844 266212
rect 429896 266200 429902 266212
rect 438854 266200 438860 266212
rect 429896 266172 438860 266200
rect 429896 266160 429902 266172
rect 438854 266160 438860 266172
rect 438912 266160 438918 266212
rect 489886 266200 489914 266240
rect 508866 266228 508872 266280
rect 508924 266268 508930 266280
rect 509142 266268 509148 266280
rect 508924 266240 509148 266268
rect 508924 266228 508930 266240
rect 509142 266228 509148 266240
rect 509200 266268 509206 266280
rect 513466 266268 513472 266280
rect 509200 266240 513472 266268
rect 509200 266228 509206 266240
rect 513466 266228 513472 266240
rect 513524 266228 513530 266280
rect 508884 266200 508912 266228
rect 489886 266172 508912 266200
rect 307018 266092 307024 266144
rect 307076 266132 307082 266144
rect 366910 266132 366916 266144
rect 307076 266104 366916 266132
rect 307076 266092 307082 266104
rect 366910 266092 366916 266104
rect 366968 266092 366974 266144
rect 360194 265684 360200 265736
rect 360252 265724 360258 265736
rect 360930 265724 360936 265736
rect 360252 265696 360936 265724
rect 360252 265684 360258 265696
rect 360930 265684 360936 265696
rect 360988 265724 360994 265736
rect 431954 265724 431960 265736
rect 360988 265696 431960 265724
rect 360988 265684 360994 265696
rect 431954 265684 431960 265696
rect 432012 265724 432018 265736
rect 432874 265724 432880 265736
rect 432012 265696 432880 265724
rect 432012 265684 432018 265696
rect 432874 265684 432880 265696
rect 432932 265724 432938 265736
rect 503714 265724 503720 265736
rect 432932 265696 503720 265724
rect 432932 265684 432938 265696
rect 503714 265684 503720 265696
rect 503772 265684 503778 265736
rect 370222 265616 370228 265668
rect 370280 265656 370286 265668
rect 440602 265656 440608 265668
rect 370280 265628 440608 265656
rect 370280 265616 370286 265628
rect 440602 265616 440608 265628
rect 440660 265656 440666 265668
rect 441062 265656 441068 265668
rect 440660 265628 441068 265656
rect 440660 265616 440666 265628
rect 441062 265616 441068 265628
rect 441120 265656 441126 265668
rect 512638 265656 512644 265668
rect 441120 265628 512644 265656
rect 441120 265616 441126 265628
rect 512638 265616 512644 265628
rect 512696 265616 512702 265668
rect 182818 264936 182824 264988
rect 182876 264976 182882 264988
rect 197354 264976 197360 264988
rect 182876 264948 197360 264976
rect 182876 264936 182882 264948
rect 197354 264936 197360 264948
rect 197412 264936 197418 264988
rect 502978 264936 502984 264988
rect 503036 264976 503042 264988
rect 510890 264976 510896 264988
rect 503036 264948 510896 264976
rect 503036 264936 503042 264948
rect 510890 264936 510896 264948
rect 510948 264936 510954 264988
rect 302694 264868 302700 264920
rect 302752 264908 302758 264920
rect 358078 264908 358084 264920
rect 302752 264880 358084 264908
rect 302752 264868 302758 264880
rect 358078 264868 358084 264880
rect 358136 264868 358142 264920
rect 302878 264188 302884 264240
rect 302936 264228 302942 264240
rect 369486 264228 369492 264240
rect 302936 264200 369492 264228
rect 302936 264188 302942 264200
rect 369486 264188 369492 264200
rect 369544 264188 369550 264240
rect 181530 262216 181536 262268
rect 181588 262256 181594 262268
rect 197354 262256 197360 262268
rect 181588 262228 197360 262256
rect 181588 262216 181594 262228
rect 197354 262216 197360 262228
rect 197412 262216 197418 262268
rect 302326 262148 302332 262200
rect 302384 262188 302390 262200
rect 359458 262188 359464 262200
rect 302384 262160 359464 262188
rect 302384 262148 302390 262160
rect 359458 262148 359464 262160
rect 359516 262148 359522 262200
rect 180150 260856 180156 260908
rect 180208 260896 180214 260908
rect 197354 260896 197360 260908
rect 180208 260868 197360 260896
rect 180208 260856 180214 260868
rect 197354 260856 197360 260868
rect 197412 260856 197418 260908
rect 357342 260108 357348 260160
rect 357400 260148 357406 260160
rect 370498 260148 370504 260160
rect 357400 260120 370504 260148
rect 357400 260108 357406 260120
rect 370498 260108 370504 260120
rect 370556 260108 370562 260160
rect 313182 258680 313188 258732
rect 313240 258720 313246 258732
rect 347682 258720 347688 258732
rect 313240 258692 347688 258720
rect 313240 258680 313246 258692
rect 347682 258680 347688 258692
rect 347740 258720 347746 258732
rect 442074 258720 442080 258732
rect 347740 258692 442080 258720
rect 347740 258680 347746 258692
rect 442074 258680 442080 258692
rect 442132 258680 442138 258732
rect 178770 258068 178776 258120
rect 178828 258108 178834 258120
rect 197354 258108 197360 258120
rect 178828 258080 197360 258108
rect 178828 258068 178834 258080
rect 197354 258068 197360 258080
rect 197412 258068 197418 258120
rect 302602 258068 302608 258120
rect 302660 258108 302666 258120
rect 313182 258108 313188 258120
rect 302660 258080 313188 258108
rect 302660 258068 302666 258080
rect 313182 258068 313188 258080
rect 313240 258068 313246 258120
rect 196618 256708 196624 256760
rect 196676 256748 196682 256760
rect 198366 256748 198372 256760
rect 196676 256720 198372 256748
rect 196676 256708 196682 256720
rect 198366 256708 198372 256720
rect 198424 256708 198430 256760
rect 302786 255960 302792 256012
rect 302844 256000 302850 256012
rect 357342 256000 357348 256012
rect 302844 255972 357348 256000
rect 302844 255960 302850 255972
rect 357342 255960 357348 255972
rect 357400 255960 357406 256012
rect 357342 255280 357348 255332
rect 357400 255320 357406 255332
rect 441706 255320 441712 255332
rect 357400 255292 441712 255320
rect 357400 255280 357406 255292
rect 441706 255280 441712 255292
rect 441764 255280 441770 255332
rect 195238 253920 195244 253972
rect 195296 253960 195302 253972
rect 197998 253960 198004 253972
rect 195296 253932 198004 253960
rect 195296 253920 195302 253932
rect 197998 253920 198004 253932
rect 198056 253920 198062 253972
rect 192570 251200 192576 251252
rect 192628 251240 192634 251252
rect 197906 251240 197912 251252
rect 192628 251212 197912 251240
rect 192628 251200 192634 251212
rect 197906 251200 197912 251212
rect 197964 251200 197970 251252
rect 302970 251200 302976 251252
rect 303028 251240 303034 251252
rect 307662 251240 307668 251252
rect 303028 251212 307668 251240
rect 303028 251200 303034 251212
rect 307662 251200 307668 251212
rect 307720 251240 307726 251252
rect 441798 251240 441804 251252
rect 307720 251212 441804 251240
rect 307720 251200 307726 251212
rect 441798 251200 441804 251212
rect 441856 251200 441862 251252
rect 303338 250452 303344 250504
rect 303396 250492 303402 250504
rect 370406 250492 370412 250504
rect 303396 250464 370412 250492
rect 303396 250452 303402 250464
rect 370406 250452 370412 250464
rect 370464 250452 370470 250504
rect 191190 249772 191196 249824
rect 191248 249812 191254 249824
rect 198090 249812 198096 249824
rect 191248 249784 198096 249812
rect 191248 249772 191254 249784
rect 198090 249772 198096 249784
rect 198148 249772 198154 249824
rect 370406 249024 370412 249076
rect 370464 249064 370470 249076
rect 388438 249064 388444 249076
rect 370464 249036 388444 249064
rect 370464 249024 370470 249036
rect 388438 249024 388444 249036
rect 388496 249064 388502 249076
rect 441890 249064 441896 249076
rect 388496 249036 441896 249064
rect 388496 249024 388502 249036
rect 441890 249024 441896 249036
rect 441948 249024 441954 249076
rect 302786 248412 302792 248464
rect 302844 248452 302850 248464
rect 370406 248452 370412 248464
rect 302844 248424 370412 248452
rect 302844 248412 302850 248424
rect 370406 248412 370412 248424
rect 370464 248412 370470 248464
rect 444374 247868 444380 247920
rect 444432 247908 444438 247920
rect 445202 247908 445208 247920
rect 444432 247880 445208 247908
rect 444432 247868 444438 247880
rect 445202 247868 445208 247880
rect 445260 247868 445266 247920
rect 371050 247664 371056 247716
rect 371108 247704 371114 247716
rect 444374 247704 444380 247716
rect 371108 247676 444380 247704
rect 371108 247664 371114 247676
rect 444374 247664 444380 247676
rect 444432 247664 444438 247716
rect 446674 247664 446680 247716
rect 446732 247704 446738 247716
rect 521930 247704 521936 247716
rect 446732 247676 521936 247704
rect 446732 247664 446738 247676
rect 521930 247664 521936 247676
rect 521988 247664 521994 247716
rect 177390 247052 177396 247104
rect 177448 247092 177454 247104
rect 197538 247092 197544 247104
rect 177448 247064 197544 247092
rect 177448 247052 177454 247064
rect 197538 247052 197544 247064
rect 197596 247052 197602 247104
rect 370498 247052 370504 247104
rect 370556 247092 370562 247104
rect 371050 247092 371056 247104
rect 370556 247064 371056 247092
rect 370556 247052 370562 247064
rect 371050 247052 371056 247064
rect 371108 247052 371114 247104
rect 340322 246304 340328 246356
rect 340380 246344 340386 246356
rect 400858 246344 400864 246356
rect 340380 246316 400864 246344
rect 340380 246304 340386 246316
rect 400858 246304 400864 246316
rect 400916 246344 400922 246356
rect 441982 246344 441988 246356
rect 400916 246316 441988 246344
rect 400916 246304 400922 246316
rect 441982 246304 441988 246316
rect 442040 246304 442046 246356
rect 302510 245624 302516 245676
rect 302568 245664 302574 245676
rect 340322 245664 340328 245676
rect 302568 245636 340328 245664
rect 302568 245624 302574 245636
rect 340322 245624 340328 245636
rect 340380 245664 340386 245676
rect 340782 245664 340788 245676
rect 340380 245636 340788 245664
rect 340380 245624 340386 245636
rect 340782 245624 340788 245636
rect 340840 245624 340846 245676
rect 312538 245556 312544 245608
rect 312596 245596 312602 245608
rect 580166 245596 580172 245608
rect 312596 245568 580172 245596
rect 312596 245556 312602 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 446490 243516 446496 243568
rect 446548 243556 446554 243568
rect 446858 243556 446864 243568
rect 446548 243528 446864 243556
rect 446548 243516 446554 243528
rect 446858 243516 446864 243528
rect 446916 243556 446922 243568
rect 517790 243556 517796 243568
rect 446916 243528 517796 243556
rect 446916 243516 446922 243528
rect 517790 243516 517796 243528
rect 517848 243556 517854 243568
rect 517974 243556 517980 243568
rect 517848 243528 517980 243556
rect 517848 243516 517854 243528
rect 517974 243516 517980 243528
rect 518032 243516 518038 243568
rect 171778 242904 171784 242956
rect 171836 242944 171842 242956
rect 197538 242944 197544 242956
rect 171836 242916 197544 242944
rect 171836 242904 171842 242916
rect 197538 242904 197544 242916
rect 197596 242904 197602 242956
rect 303246 242904 303252 242956
rect 303304 242944 303310 242956
rect 443546 242944 443552 242956
rect 303304 242916 443552 242944
rect 303304 242904 303310 242916
rect 443546 242904 443552 242916
rect 443604 242904 443610 242956
rect 377398 242836 377404 242888
rect 377456 242876 377462 242888
rect 377766 242876 377772 242888
rect 377456 242848 377772 242876
rect 377456 242836 377462 242848
rect 377766 242836 377772 242848
rect 377824 242876 377830 242888
rect 444466 242876 444472 242888
rect 377824 242848 444472 242876
rect 377824 242836 377830 242848
rect 444466 242836 444472 242848
rect 444524 242876 444530 242888
rect 444926 242876 444932 242888
rect 444524 242848 444932 242876
rect 444524 242836 444530 242848
rect 444926 242836 444932 242848
rect 444984 242836 444990 242888
rect 342898 242156 342904 242208
rect 342956 242196 342962 242208
rect 377766 242196 377772 242208
rect 342956 242168 377772 242196
rect 342956 242156 342962 242168
rect 377766 242156 377772 242168
rect 377824 242156 377830 242208
rect 195330 241476 195336 241528
rect 195388 241516 195394 241528
rect 198274 241516 198280 241528
rect 195388 241488 198280 241516
rect 195388 241476 195394 241488
rect 198274 241476 198280 241488
rect 198332 241476 198338 241528
rect 444558 241408 444564 241460
rect 444616 241448 444622 241460
rect 444834 241448 444840 241460
rect 444616 241420 444840 241448
rect 444616 241408 444622 241420
rect 444834 241408 444840 241420
rect 444892 241408 444898 241460
rect 446490 241408 446496 241460
rect 446548 241448 446554 241460
rect 446766 241448 446772 241460
rect 446548 241420 446772 241448
rect 446548 241408 446554 241420
rect 446766 241408 446772 241420
rect 446824 241408 446830 241460
rect 304258 240728 304264 240780
rect 304316 240768 304322 240780
rect 374546 240768 374552 240780
rect 304316 240740 374552 240768
rect 304316 240728 304322 240740
rect 374546 240728 374552 240740
rect 374604 240768 374610 240780
rect 406378 240768 406384 240780
rect 374604 240740 406384 240768
rect 374604 240728 374610 240740
rect 406378 240728 406384 240740
rect 406436 240728 406442 240780
rect 446490 240728 446496 240780
rect 446548 240768 446554 240780
rect 519170 240768 519176 240780
rect 446548 240740 519176 240768
rect 446548 240728 446554 240740
rect 519170 240728 519176 240740
rect 519228 240728 519234 240780
rect 406378 240116 406384 240168
rect 406436 240156 406442 240168
rect 444558 240156 444564 240168
rect 406436 240128 444564 240156
rect 406436 240116 406442 240128
rect 444558 240116 444564 240128
rect 444616 240116 444622 240168
rect 444650 240048 444656 240100
rect 444708 240088 444714 240100
rect 445202 240088 445208 240100
rect 444708 240060 445208 240088
rect 444708 240048 444714 240060
rect 445202 240048 445208 240060
rect 445260 240048 445266 240100
rect 445202 239368 445208 239420
rect 445260 239408 445266 239420
rect 517882 239408 517888 239420
rect 445260 239380 517888 239408
rect 445260 239368 445266 239380
rect 517882 239368 517888 239380
rect 517940 239368 517946 239420
rect 171870 238756 171876 238808
rect 171928 238796 171934 238808
rect 197538 238796 197544 238808
rect 171928 238768 197544 238796
rect 171928 238756 171934 238768
rect 197538 238756 197544 238768
rect 197596 238756 197602 238808
rect 443638 238348 443644 238400
rect 443696 238388 443702 238400
rect 444282 238388 444288 238400
rect 443696 238360 444288 238388
rect 443696 238348 443702 238360
rect 444282 238348 444288 238360
rect 444340 238348 444346 238400
rect 444282 238008 444288 238060
rect 444340 238048 444346 238060
rect 523126 238048 523132 238060
rect 444340 238020 523132 238048
rect 444340 238008 444346 238020
rect 523126 238008 523132 238020
rect 523184 238008 523190 238060
rect 196710 237736 196716 237788
rect 196768 237776 196774 237788
rect 198458 237776 198464 237788
rect 196768 237748 198464 237776
rect 196768 237736 196774 237748
rect 198458 237736 198464 237748
rect 198516 237736 198522 237788
rect 378226 236648 378232 236700
rect 378284 236688 378290 236700
rect 443178 236688 443184 236700
rect 378284 236660 443184 236688
rect 378284 236648 378290 236660
rect 443178 236648 443184 236660
rect 443236 236648 443242 236700
rect 446582 236648 446588 236700
rect 446640 236688 446646 236700
rect 519078 236688 519084 236700
rect 446640 236660 519084 236688
rect 446640 236648 446646 236660
rect 519078 236648 519084 236660
rect 519136 236648 519142 236700
rect 302786 235968 302792 236020
rect 302844 236008 302850 236020
rect 375466 236008 375472 236020
rect 302844 235980 375472 236008
rect 302844 235968 302850 235980
rect 375466 235968 375472 235980
rect 375524 236008 375530 236020
rect 378226 236008 378232 236020
rect 375524 235980 378232 236008
rect 375524 235968 375530 235980
rect 378226 235968 378232 235980
rect 378284 235968 378290 236020
rect 447962 235220 447968 235272
rect 448020 235260 448026 235272
rect 521746 235260 521752 235272
rect 448020 235232 521752 235260
rect 448020 235220 448026 235232
rect 521746 235220 521752 235232
rect 521804 235260 521810 235272
rect 522022 235260 522028 235272
rect 521804 235232 522028 235260
rect 521804 235220 521810 235232
rect 522022 235220 522028 235232
rect 522080 235220 522086 235272
rect 171962 234608 171968 234660
rect 172020 234648 172026 234660
rect 197538 234648 197544 234660
rect 172020 234620 197544 234648
rect 172020 234608 172026 234620
rect 197538 234608 197544 234620
rect 197596 234608 197602 234660
rect 516226 234540 516232 234592
rect 516284 234580 516290 234592
rect 518894 234580 518900 234592
rect 516284 234552 518900 234580
rect 516284 234540 516290 234552
rect 518894 234540 518900 234552
rect 518952 234540 518958 234592
rect 376662 233860 376668 233912
rect 376720 233900 376726 233912
rect 385678 233900 385684 233912
rect 376720 233872 385684 233900
rect 376720 233860 376726 233872
rect 385678 233860 385684 233872
rect 385736 233900 385742 233912
rect 443270 233900 443276 233912
rect 385736 233872 443276 233900
rect 385736 233860 385742 233872
rect 443270 233860 443276 233872
rect 443328 233860 443334 233912
rect 445294 233860 445300 233912
rect 445352 233900 445358 233912
rect 528646 233900 528652 233912
rect 445352 233872 528652 233900
rect 445352 233860 445358 233872
rect 528646 233860 528652 233872
rect 528704 233860 528710 233912
rect 172054 233248 172060 233300
rect 172112 233288 172118 233300
rect 197354 233288 197360 233300
rect 172112 233260 197360 233288
rect 172112 233248 172118 233260
rect 197354 233248 197360 233260
rect 197412 233248 197418 233300
rect 302694 233248 302700 233300
rect 302752 233288 302758 233300
rect 375558 233288 375564 233300
rect 302752 233260 375564 233288
rect 302752 233248 302758 233260
rect 375558 233248 375564 233260
rect 375616 233288 375622 233300
rect 376662 233288 376668 233300
rect 375616 233260 376668 233288
rect 375616 233248 375622 233260
rect 376662 233248 376668 233260
rect 376720 233248 376726 233300
rect 449250 233248 449256 233300
rect 449308 233288 449314 233300
rect 516226 233288 516232 233300
rect 449308 233260 516232 233288
rect 449308 233248 449314 233260
rect 516226 233248 516232 233260
rect 516284 233288 516290 233300
rect 516594 233288 516600 233300
rect 516284 233260 516600 233288
rect 516284 233248 516290 233260
rect 516594 233248 516600 233260
rect 516652 233248 516658 233300
rect 447870 233180 447876 233232
rect 447928 233220 447934 233232
rect 448146 233220 448152 233232
rect 447928 233192 448152 233220
rect 447928 233180 447934 233192
rect 448146 233180 448152 233192
rect 448204 233180 448210 233232
rect 516410 233180 516416 233232
rect 516468 233220 516474 233232
rect 519262 233220 519268 233232
rect 516468 233192 519268 233220
rect 516468 233180 516474 233192
rect 519262 233180 519268 233192
rect 519320 233180 519326 233232
rect 448146 231820 448152 231872
rect 448204 231860 448210 231872
rect 516410 231860 516416 231872
rect 448204 231832 516416 231860
rect 448204 231820 448210 231832
rect 516410 231820 516416 231832
rect 516468 231820 516474 231872
rect 375650 231072 375656 231124
rect 375708 231112 375714 231124
rect 380894 231112 380900 231124
rect 375708 231084 380900 231112
rect 375708 231072 375714 231084
rect 380894 231072 380900 231084
rect 380952 231112 380958 231124
rect 443362 231112 443368 231124
rect 380952 231084 443368 231112
rect 380952 231072 380958 231084
rect 443362 231072 443368 231084
rect 443420 231072 443426 231124
rect 444926 231072 444932 231124
rect 444984 231112 444990 231124
rect 521838 231112 521844 231124
rect 444984 231084 521844 231112
rect 444984 231072 444990 231084
rect 521838 231072 521844 231084
rect 521896 231072 521902 231124
rect 302786 230460 302792 230512
rect 302844 230500 302850 230512
rect 375650 230500 375656 230512
rect 302844 230472 375656 230500
rect 302844 230460 302850 230472
rect 375650 230460 375656 230472
rect 375708 230460 375714 230512
rect 444834 230392 444840 230444
rect 444892 230432 444898 230444
rect 445110 230432 445116 230444
rect 444892 230404 445116 230432
rect 444892 230392 444898 230404
rect 445110 230392 445116 230404
rect 445168 230392 445174 230444
rect 371142 229712 371148 229764
rect 371200 229752 371206 229764
rect 444834 229752 444840 229764
rect 371200 229724 444840 229752
rect 371200 229712 371206 229724
rect 444834 229712 444840 229724
rect 444892 229712 444898 229764
rect 446398 229712 446404 229764
rect 446456 229752 446462 229764
rect 520550 229752 520556 229764
rect 446456 229724 520556 229752
rect 446456 229712 446462 229724
rect 520550 229712 520556 229724
rect 520608 229712 520614 229764
rect 174630 229100 174636 229152
rect 174688 229140 174694 229152
rect 197354 229140 197360 229152
rect 174688 229112 197360 229140
rect 174688 229100 174694 229112
rect 197354 229100 197360 229112
rect 197412 229100 197418 229152
rect 517698 228692 517704 228744
rect 517756 228732 517762 228744
rect 518250 228732 518256 228744
rect 517756 228704 518256 228732
rect 517756 228692 517762 228704
rect 518250 228692 518256 228704
rect 518308 228692 518314 228744
rect 448054 228420 448060 228472
rect 448112 228460 448118 228472
rect 517698 228460 517704 228472
rect 448112 228432 517704 228460
rect 448112 228420 448118 228432
rect 517698 228420 517704 228432
rect 517756 228420 517762 228472
rect 445386 228352 445392 228404
rect 445444 228392 445450 228404
rect 524598 228392 524604 228404
rect 445444 228364 524604 228392
rect 445444 228352 445450 228364
rect 524598 228352 524604 228364
rect 524656 228352 524662 228404
rect 441798 228284 441804 228336
rect 441856 228324 441862 228336
rect 442350 228324 442356 228336
rect 441856 228296 442356 228324
rect 441856 228284 441862 228296
rect 442350 228284 442356 228296
rect 442408 228284 442414 228336
rect 447870 227740 447876 227792
rect 447928 227780 447934 227792
rect 448054 227780 448060 227792
rect 447928 227752 448060 227780
rect 447928 227740 447934 227752
rect 448054 227740 448060 227752
rect 448112 227740 448118 227792
rect 302786 227672 302792 227724
rect 302844 227712 302850 227724
rect 382274 227712 382280 227724
rect 302844 227684 382280 227712
rect 302844 227672 302850 227684
rect 382274 227672 382280 227684
rect 382332 227672 382338 227724
rect 382274 226992 382280 227044
rect 382332 227032 382338 227044
rect 394142 227032 394148 227044
rect 382332 227004 394148 227032
rect 382332 226992 382338 227004
rect 394142 226992 394148 227004
rect 394200 226992 394206 227044
rect 516226 226788 516232 226840
rect 516284 226828 516290 226840
rect 520458 226828 520464 226840
rect 516284 226800 520464 226828
rect 516284 226788 516290 226800
rect 520458 226788 520464 226800
rect 520516 226788 520522 226840
rect 176010 226312 176016 226364
rect 176068 226352 176074 226364
rect 197538 226352 197544 226364
rect 176068 226324 197544 226352
rect 176068 226312 176074 226324
rect 197538 226312 197544 226324
rect 197596 226312 197602 226364
rect 394142 226312 394148 226364
rect 394200 226352 394206 226364
rect 394602 226352 394608 226364
rect 394200 226324 394608 226352
rect 394200 226312 394206 226324
rect 394602 226312 394608 226324
rect 394660 226352 394666 226364
rect 443454 226352 443460 226364
rect 394660 226324 443460 226352
rect 394660 226312 394666 226324
rect 443454 226312 443460 226324
rect 443512 226312 443518 226364
rect 447778 226312 447784 226364
rect 447836 226352 447842 226364
rect 516226 226352 516232 226364
rect 447836 226324 516232 226352
rect 447836 226312 447842 226324
rect 516226 226312 516232 226324
rect 516284 226352 516290 226364
rect 516502 226352 516508 226364
rect 516284 226324 516508 226352
rect 516284 226312 516290 226324
rect 516502 226312 516508 226324
rect 516560 226312 516566 226364
rect 375190 226244 375196 226296
rect 375248 226284 375254 226296
rect 441614 226284 441620 226296
rect 375248 226256 441620 226284
rect 375248 226244 375254 226256
rect 441614 226244 441620 226256
rect 441672 226244 441678 226296
rect 516134 226244 516140 226296
rect 516192 226284 516198 226296
rect 524506 226284 524512 226296
rect 516192 226256 524512 226284
rect 516192 226244 516198 226256
rect 524506 226244 524512 226256
rect 524564 226244 524570 226296
rect 375098 226176 375104 226228
rect 375156 226216 375162 226228
rect 375156 226188 431954 226216
rect 375156 226176 375162 226188
rect 431926 226148 431954 226188
rect 441614 226148 441620 226160
rect 431926 226120 441620 226148
rect 441614 226108 441620 226120
rect 441672 226108 441678 226160
rect 304902 225632 304908 225684
rect 304960 225672 304966 225684
rect 367830 225672 367836 225684
rect 304960 225644 367836 225672
rect 304960 225632 304966 225644
rect 367830 225632 367836 225644
rect 367888 225632 367894 225684
rect 509142 225632 509148 225684
rect 509200 225672 509206 225684
rect 514846 225672 514852 225684
rect 509200 225644 514852 225672
rect 509200 225632 509206 225644
rect 514846 225632 514852 225644
rect 514904 225632 514910 225684
rect 302970 225564 302976 225616
rect 303028 225604 303034 225616
rect 371142 225604 371148 225616
rect 303028 225576 371148 225604
rect 303028 225564 303034 225576
rect 371142 225564 371148 225576
rect 371200 225564 371206 225616
rect 507762 225564 507768 225616
rect 507820 225604 507826 225616
rect 507820 225576 509234 225604
rect 507820 225564 507826 225576
rect 509206 225536 509234 225576
rect 512638 225564 512644 225616
rect 512696 225604 512702 225616
rect 514938 225604 514944 225616
rect 512696 225576 514944 225604
rect 512696 225564 512702 225576
rect 514938 225564 514944 225576
rect 514996 225564 515002 225616
rect 514754 225536 514760 225548
rect 509206 225508 514760 225536
rect 514754 225496 514760 225508
rect 514812 225496 514818 225548
rect 441982 225156 441988 225208
rect 442040 225196 442046 225208
rect 442258 225196 442264 225208
rect 442040 225168 442264 225196
rect 442040 225156 442046 225168
rect 442258 225156 442264 225168
rect 442316 225156 442322 225208
rect 441890 225088 441896 225140
rect 441948 225128 441954 225140
rect 442166 225128 442172 225140
rect 441948 225100 442172 225128
rect 441948 225088 441954 225100
rect 442166 225088 442172 225100
rect 442224 225088 442230 225140
rect 351914 225020 351920 225072
rect 351972 225060 351978 225072
rect 375834 225060 375840 225072
rect 351972 225032 375840 225060
rect 351972 225020 351978 225032
rect 375834 225020 375840 225032
rect 375892 225060 375898 225072
rect 445938 225060 445944 225072
rect 375892 225032 445944 225060
rect 375892 225020 375898 225032
rect 445938 225020 445944 225032
rect 445996 225020 446002 225072
rect 464338 225020 464344 225072
rect 464396 225060 464402 225072
rect 513742 225060 513748 225072
rect 464396 225032 513748 225060
rect 464396 225020 464402 225032
rect 513742 225020 513748 225032
rect 513800 225020 513806 225072
rect 177298 224952 177304 225004
rect 177356 224992 177362 225004
rect 197354 224992 197360 225004
rect 177356 224964 197360 224992
rect 177356 224952 177362 224964
rect 197354 224952 197360 224964
rect 197412 224952 197418 225004
rect 345658 224952 345664 225004
rect 345716 224992 345722 225004
rect 375742 224992 375748 225004
rect 345716 224964 375748 224992
rect 345716 224952 345722 224964
rect 375742 224952 375748 224964
rect 375800 224992 375806 225004
rect 445846 224992 445852 225004
rect 375800 224964 445852 224992
rect 375800 224952 375806 224964
rect 445846 224952 445852 224964
rect 445904 224952 445910 225004
rect 456058 224952 456064 225004
rect 456116 224992 456122 225004
rect 513374 224992 513380 225004
rect 456116 224964 513380 224992
rect 456116 224952 456122 224964
rect 513374 224952 513380 224964
rect 513432 224952 513438 225004
rect 390462 224884 390468 224936
rect 390520 224924 390526 224936
rect 441706 224924 441712 224936
rect 390520 224896 441712 224924
rect 390520 224884 390526 224896
rect 441706 224884 441712 224896
rect 441764 224884 441770 224936
rect 516134 224884 516140 224936
rect 516192 224924 516198 224936
rect 521654 224924 521660 224936
rect 516192 224896 521660 224924
rect 516192 224884 516198 224896
rect 521654 224884 521660 224896
rect 521712 224884 521718 224936
rect 393222 224816 393228 224868
rect 393280 224856 393286 224868
rect 441614 224856 441620 224868
rect 393280 224828 441620 224856
rect 393280 224816 393286 224828
rect 441614 224816 441620 224828
rect 441672 224816 441678 224868
rect 302878 224340 302884 224392
rect 302936 224380 302942 224392
rect 340874 224380 340880 224392
rect 302936 224352 340880 224380
rect 302936 224340 302942 224352
rect 340874 224340 340880 224352
rect 340932 224340 340938 224392
rect 358078 224272 358084 224324
rect 358136 224312 358142 224324
rect 369394 224312 369400 224324
rect 358136 224284 369400 224312
rect 358136 224272 358142 224284
rect 369394 224272 369400 224284
rect 369452 224312 369458 224324
rect 371326 224312 371332 224324
rect 369452 224284 371332 224312
rect 369452 224272 369458 224284
rect 371326 224272 371332 224284
rect 371384 224272 371390 224324
rect 444466 224272 444472 224324
rect 444524 224312 444530 224324
rect 445570 224312 445576 224324
rect 444524 224284 445576 224312
rect 444524 224272 444530 224284
rect 445570 224272 445576 224284
rect 445628 224272 445634 224324
rect 302878 224204 302884 224256
rect 302936 224244 302942 224256
rect 370498 224244 370504 224256
rect 302936 224216 370504 224244
rect 302936 224204 302942 224216
rect 370498 224204 370504 224216
rect 370556 224204 370562 224256
rect 378134 224204 378140 224256
rect 378192 224244 378198 224256
rect 443178 224244 443184 224256
rect 378192 224216 443184 224244
rect 378192 224204 378198 224216
rect 443178 224204 443184 224216
rect 443236 224204 443242 224256
rect 445110 224204 445116 224256
rect 445168 224244 445174 224256
rect 445662 224244 445668 224256
rect 445168 224216 445668 224244
rect 445168 224204 445174 224216
rect 445662 224204 445668 224216
rect 445720 224204 445726 224256
rect 302326 223932 302332 223984
rect 302384 223972 302390 223984
rect 375926 223972 375932 223984
rect 302384 223944 375932 223972
rect 302384 223932 302390 223944
rect 375926 223932 375932 223944
rect 375984 223972 375990 223984
rect 378134 223972 378140 223984
rect 375984 223944 378140 223972
rect 375984 223932 375990 223944
rect 378134 223932 378140 223944
rect 378192 223932 378198 223984
rect 340874 223864 340880 223916
rect 340932 223904 340938 223916
rect 342162 223904 342168 223916
rect 340932 223876 342168 223904
rect 340932 223864 340938 223876
rect 342162 223864 342168 223876
rect 342220 223904 342226 223916
rect 441798 223904 441804 223916
rect 342220 223876 441804 223904
rect 342220 223864 342226 223876
rect 441798 223864 441804 223876
rect 441856 223864 441862 223916
rect 461578 223864 461584 223916
rect 461636 223904 461642 223916
rect 513742 223904 513748 223916
rect 461636 223876 513748 223904
rect 461636 223864 461642 223876
rect 513742 223864 513748 223876
rect 513800 223864 513806 223916
rect 170490 222844 170496 222896
rect 170548 222884 170554 222896
rect 198182 222884 198188 222896
rect 170548 222856 198188 222884
rect 170548 222844 170554 222856
rect 198182 222844 198188 222856
rect 198240 222844 198246 222896
rect 444742 222300 444748 222352
rect 444800 222340 444806 222352
rect 483658 222340 483664 222352
rect 444800 222312 483664 222340
rect 444800 222300 444806 222312
rect 483658 222300 483664 222312
rect 483716 222300 483722 222352
rect 445570 222232 445576 222284
rect 445628 222272 445634 222284
rect 489178 222272 489184 222284
rect 445628 222244 489184 222272
rect 445628 222232 445634 222244
rect 489178 222232 489184 222244
rect 489236 222232 489242 222284
rect 445662 222164 445668 222216
rect 445720 222204 445726 222216
rect 485038 222204 485044 222216
rect 445720 222176 485044 222204
rect 445720 222164 445726 222176
rect 485038 222164 485044 222176
rect 485096 222164 485102 222216
rect 302326 222096 302332 222148
rect 302384 222136 302390 222148
rect 351914 222136 351920 222148
rect 302384 222108 351920 222136
rect 302384 222096 302390 222108
rect 351914 222096 351920 222108
rect 351972 222096 351978 222148
rect 454678 222096 454684 222148
rect 454736 222136 454742 222148
rect 456058 222136 456064 222148
rect 454736 222108 456064 222136
rect 454736 222096 454742 222108
rect 456058 222096 456064 222108
rect 456116 222096 456122 222148
rect 516134 222096 516140 222148
rect 516192 222136 516198 222148
rect 524414 222136 524420 222148
rect 516192 222108 524420 222136
rect 516192 222096 516198 222108
rect 524414 222096 524420 222108
rect 524472 222096 524478 222148
rect 191098 220872 191104 220924
rect 191156 220912 191162 220924
rect 197354 220912 197360 220924
rect 191156 220884 197360 220912
rect 191156 220872 191162 220884
rect 197354 220872 197360 220884
rect 197412 220872 197418 220924
rect 370314 220872 370320 220924
rect 370372 220912 370378 220924
rect 376018 220912 376024 220924
rect 370372 220884 376024 220912
rect 370372 220872 370378 220884
rect 376018 220872 376024 220884
rect 376076 220872 376082 220924
rect 444742 220872 444748 220924
rect 444800 220912 444806 220924
rect 482278 220912 482284 220924
rect 444800 220884 482284 220912
rect 444800 220872 444806 220884
rect 482278 220872 482284 220884
rect 482336 220872 482342 220924
rect 445570 220804 445576 220856
rect 445628 220844 445634 220856
rect 490558 220844 490564 220856
rect 445628 220816 490564 220844
rect 445628 220804 445634 220816
rect 490558 220804 490564 220816
rect 490616 220804 490622 220856
rect 371510 220736 371516 220788
rect 371568 220776 371574 220788
rect 372430 220776 372436 220788
rect 371568 220748 372436 220776
rect 371568 220736 371574 220748
rect 372430 220736 372436 220748
rect 372488 220776 372494 220788
rect 376110 220776 376116 220788
rect 372488 220748 376116 220776
rect 372488 220736 372494 220748
rect 376110 220736 376116 220748
rect 376168 220736 376174 220788
rect 516134 220736 516140 220788
rect 516192 220776 516198 220788
rect 523126 220776 523132 220788
rect 516192 220748 523132 220776
rect 516192 220736 516198 220748
rect 523126 220736 523132 220748
rect 523184 220736 523190 220788
rect 516134 219920 516140 219972
rect 516192 219960 516198 219972
rect 517974 219960 517980 219972
rect 516192 219932 517980 219960
rect 516192 219920 516198 219932
rect 517974 219920 517980 219932
rect 518032 219920 518038 219972
rect 445662 219580 445668 219632
rect 445720 219620 445726 219632
rect 479518 219620 479524 219632
rect 445720 219592 479524 219620
rect 445720 219580 445726 219592
rect 479518 219580 479524 219592
rect 479576 219580 479582 219632
rect 443270 219512 443276 219564
rect 443328 219512 443334 219564
rect 444742 219512 444748 219564
rect 444800 219552 444806 219564
rect 493318 219552 493324 219564
rect 444800 219524 493324 219552
rect 444800 219512 444806 219524
rect 493318 219512 493324 219524
rect 493376 219512 493382 219564
rect 302418 219376 302424 219428
rect 302476 219416 302482 219428
rect 345658 219416 345664 219428
rect 302476 219388 345664 219416
rect 302476 219376 302482 219388
rect 345658 219376 345664 219388
rect 345716 219376 345722 219428
rect 443288 219416 443316 219512
rect 445570 219444 445576 219496
rect 445628 219484 445634 219496
rect 494698 219484 494704 219496
rect 445628 219456 494704 219484
rect 445628 219444 445634 219456
rect 494698 219444 494704 219456
rect 494756 219444 494762 219496
rect 443638 219416 443644 219428
rect 443288 219388 443644 219416
rect 443638 219376 443644 219388
rect 443696 219376 443702 219428
rect 519538 219376 519544 219428
rect 519596 219416 519602 219428
rect 580166 219416 580172 219428
rect 519596 219388 580172 219416
rect 519596 219376 519602 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 516134 219308 516140 219360
rect 516192 219348 516198 219360
rect 522022 219348 522028 219360
rect 516192 219320 522028 219348
rect 516192 219308 516198 219320
rect 522022 219308 522028 219320
rect 522080 219308 522086 219360
rect 370314 218424 370320 218476
rect 370372 218464 370378 218476
rect 374178 218464 374184 218476
rect 370372 218436 374184 218464
rect 370372 218424 370378 218436
rect 374178 218424 374184 218436
rect 374236 218464 374242 218476
rect 374822 218464 374828 218476
rect 374236 218436 374828 218464
rect 374236 218424 374242 218436
rect 374822 218424 374828 218436
rect 374880 218424 374886 218476
rect 443638 218084 443644 218136
rect 443696 218124 443702 218136
rect 475378 218124 475384 218136
rect 443696 218096 475384 218124
rect 443696 218084 443702 218096
rect 475378 218084 475384 218096
rect 475436 218084 475442 218136
rect 192478 218016 192484 218068
rect 192536 218056 192542 218068
rect 197538 218056 197544 218068
rect 192536 218028 197544 218056
rect 192536 218016 192542 218028
rect 197538 218016 197544 218028
rect 197596 218016 197602 218068
rect 443362 218016 443368 218068
rect 443420 218056 443426 218068
rect 497458 218056 497464 218068
rect 443420 218028 497464 218056
rect 443420 218016 443426 218028
rect 497458 218016 497464 218028
rect 497516 218016 497522 218068
rect 370958 217336 370964 217388
rect 371016 217376 371022 217388
rect 372982 217376 372988 217388
rect 371016 217348 372988 217376
rect 371016 217336 371022 217348
rect 372982 217336 372988 217348
rect 373040 217336 373046 217388
rect 517054 217336 517060 217388
rect 517112 217376 517118 217388
rect 518894 217376 518900 217388
rect 517112 217348 518900 217376
rect 517112 217336 517118 217348
rect 518894 217336 518900 217348
rect 518952 217336 518958 217388
rect 445938 217268 445944 217320
rect 445996 217308 446002 217320
rect 471238 217308 471244 217320
rect 445996 217280 471244 217308
rect 445996 217268 446002 217280
rect 471238 217268 471244 217280
rect 471296 217268 471302 217320
rect 188430 216656 188436 216708
rect 188488 216696 188494 216708
rect 197354 216696 197360 216708
rect 188488 216668 197360 216696
rect 188488 216656 188494 216668
rect 197354 216656 197360 216668
rect 197412 216656 197418 216708
rect 372982 216656 372988 216708
rect 373040 216696 373046 216708
rect 373534 216696 373540 216708
rect 373040 216668 373540 216696
rect 373040 216656 373046 216668
rect 373534 216656 373540 216668
rect 373592 216656 373598 216708
rect 443270 216656 443276 216708
rect 443328 216696 443334 216708
rect 472618 216696 472624 216708
rect 443328 216668 472624 216696
rect 443328 216656 443334 216668
rect 472618 216656 472624 216668
rect 472676 216656 472682 216708
rect 516134 216588 516140 216640
rect 516192 216628 516198 216640
rect 521930 216628 521936 216640
rect 516192 216600 521936 216628
rect 516192 216588 516198 216600
rect 521930 216588 521936 216600
rect 521988 216588 521994 216640
rect 370958 216180 370964 216232
rect 371016 216220 371022 216232
rect 374638 216220 374644 216232
rect 371016 216192 374644 216220
rect 371016 216180 371022 216192
rect 374638 216180 374644 216192
rect 374696 216180 374702 216232
rect 303062 215908 303068 215960
rect 303120 215948 303126 215960
rect 303522 215948 303528 215960
rect 303120 215920 303528 215948
rect 303120 215908 303126 215920
rect 303522 215908 303528 215920
rect 303580 215948 303586 215960
rect 352558 215948 352564 215960
rect 303580 215920 352564 215948
rect 303580 215908 303586 215920
rect 352558 215908 352564 215920
rect 352616 215908 352622 215960
rect 445846 215908 445852 215960
rect 445904 215948 445910 215960
rect 468478 215948 468484 215960
rect 445904 215920 468484 215948
rect 445904 215908 445910 215920
rect 468478 215908 468484 215920
rect 468536 215908 468542 215960
rect 444466 215840 444472 215892
rect 444524 215880 444530 215892
rect 446030 215880 446036 215892
rect 444524 215852 446036 215880
rect 444524 215840 444530 215852
rect 446030 215840 446036 215852
rect 446088 215840 446094 215892
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 199378 215268 199384 215280
rect 3384 215240 199384 215268
rect 3384 215228 3390 215240
rect 199378 215228 199384 215240
rect 199436 215228 199442 215280
rect 370682 215024 370688 215076
rect 370740 215064 370746 215076
rect 374362 215064 374368 215076
rect 370740 215036 374368 215064
rect 370740 215024 370746 215036
rect 374362 215024 374368 215036
rect 374420 215024 374426 215076
rect 187050 213936 187056 213988
rect 187108 213976 187114 213988
rect 197354 213976 197360 213988
rect 187108 213948 197360 213976
rect 187108 213936 187114 213948
rect 197354 213936 197360 213948
rect 197412 213936 197418 213988
rect 372798 213868 372804 213920
rect 372856 213908 372862 213920
rect 373350 213908 373356 213920
rect 372856 213880 373356 213908
rect 372856 213868 372862 213880
rect 373350 213868 373356 213880
rect 373408 213868 373414 213920
rect 516226 213868 516232 213920
rect 516284 213908 516290 213920
rect 518066 213908 518072 213920
rect 516284 213880 518072 213908
rect 516284 213868 516290 213880
rect 518066 213868 518072 213880
rect 518124 213868 518130 213920
rect 370958 213800 370964 213852
rect 371016 213840 371022 213852
rect 374270 213840 374276 213852
rect 371016 213812 374276 213840
rect 371016 213800 371022 213812
rect 374270 213800 374276 213812
rect 374328 213800 374334 213852
rect 516134 213800 516140 213852
rect 516192 213840 516198 213852
rect 520550 213840 520556 213852
rect 516192 213812 520556 213840
rect 516192 213800 516198 213812
rect 520550 213800 520556 213812
rect 520608 213800 520614 213852
rect 445110 212848 445116 212900
rect 445168 212888 445174 212900
rect 445938 212888 445944 212900
rect 445168 212860 445944 212888
rect 445168 212848 445174 212860
rect 445938 212848 445944 212860
rect 445996 212848 446002 212900
rect 444742 212440 444748 212492
rect 444800 212480 444806 212492
rect 486418 212480 486424 212492
rect 444800 212452 486424 212480
rect 444800 212440 444806 212452
rect 486418 212440 486424 212452
rect 486476 212440 486482 212492
rect 442718 212372 442724 212424
rect 442776 212412 442782 212424
rect 445018 212412 445024 212424
rect 442776 212384 445024 212412
rect 442776 212372 442782 212384
rect 445018 212372 445024 212384
rect 445076 212412 445082 212424
rect 476758 212412 476764 212424
rect 445076 212384 476764 212412
rect 445076 212372 445082 212384
rect 476758 212372 476764 212384
rect 476816 212372 476822 212424
rect 445110 212304 445116 212356
rect 445168 212344 445174 212356
rect 457438 212344 457444 212356
rect 445168 212316 457444 212344
rect 445168 212304 445174 212316
rect 457438 212304 457444 212316
rect 457496 212304 457502 212356
rect 516134 211896 516140 211948
rect 516192 211936 516198 211948
rect 519078 211936 519084 211948
rect 516192 211908 519084 211936
rect 516192 211896 516198 211908
rect 519078 211896 519084 211908
rect 519136 211896 519142 211948
rect 370958 211556 370964 211608
rect 371016 211596 371022 211608
rect 373442 211596 373448 211608
rect 371016 211568 373448 211596
rect 371016 211556 371022 211568
rect 373442 211556 373448 211568
rect 373500 211556 373506 211608
rect 184290 211148 184296 211200
rect 184348 211188 184354 211200
rect 197354 211188 197360 211200
rect 184348 211160 197360 211188
rect 184348 211148 184354 211160
rect 197354 211148 197360 211160
rect 197412 211148 197418 211200
rect 443178 211080 443184 211132
rect 443236 211120 443242 211132
rect 448514 211120 448520 211132
rect 443236 211092 448520 211120
rect 443236 211080 443242 211092
rect 448514 211080 448520 211092
rect 448572 211080 448578 211132
rect 516410 211080 516416 211132
rect 516468 211120 516474 211132
rect 518342 211120 518348 211132
rect 516468 211092 518348 211120
rect 516468 211080 516474 211092
rect 518342 211080 518348 211092
rect 518400 211080 518406 211132
rect 442166 211012 442172 211064
rect 442224 211052 442230 211064
rect 449158 211052 449164 211064
rect 442224 211024 449164 211052
rect 442224 211012 442230 211024
rect 449158 211012 449164 211024
rect 449216 211012 449222 211064
rect 370958 210264 370964 210316
rect 371016 210304 371022 210316
rect 372706 210304 372712 210316
rect 371016 210276 372712 210304
rect 371016 210264 371022 210276
rect 372706 210264 372712 210276
rect 372764 210304 372770 210316
rect 373258 210304 373264 210316
rect 372764 210276 373264 210304
rect 372764 210264 372770 210276
rect 373258 210264 373264 210276
rect 373316 210264 373322 210316
rect 182910 209788 182916 209840
rect 182968 209828 182974 209840
rect 197354 209828 197360 209840
rect 182968 209800 197360 209828
rect 182968 209788 182974 209800
rect 197354 209788 197360 209800
rect 197412 209788 197418 209840
rect 516134 209516 516140 209568
rect 516192 209556 516198 209568
rect 519170 209556 519176 209568
rect 516192 209528 519176 209556
rect 516192 209516 516198 209528
rect 519170 209516 519176 209528
rect 519228 209516 519234 209568
rect 370958 209176 370964 209228
rect 371016 209216 371022 209228
rect 372890 209216 372896 209228
rect 371016 209188 372896 209216
rect 371016 209176 371022 209188
rect 372890 209176 372896 209188
rect 372948 209176 372954 209228
rect 445662 209108 445668 209160
rect 445720 209148 445726 209160
rect 450538 209148 450544 209160
rect 445720 209120 450544 209148
rect 445720 209108 445726 209120
rect 450538 209108 450544 209120
rect 450596 209148 450602 209160
rect 461578 209148 461584 209160
rect 450596 209120 461584 209148
rect 450596 209108 450602 209120
rect 461578 209108 461584 209120
rect 461636 209108 461642 209160
rect 303062 209040 303068 209092
rect 303120 209080 303126 209092
rect 303522 209080 303528 209092
rect 303120 209052 303528 209080
rect 303120 209040 303126 209052
rect 303522 209040 303528 209052
rect 303580 209080 303586 209092
rect 342898 209080 342904 209092
rect 303580 209052 342904 209080
rect 303580 209040 303586 209052
rect 342898 209040 342904 209052
rect 342956 209040 342962 209092
rect 444558 209040 444564 209092
rect 444616 209080 444622 209092
rect 445110 209080 445116 209092
rect 444616 209052 445116 209080
rect 444616 209040 444622 209052
rect 445110 209040 445116 209052
rect 445168 209080 445174 209092
rect 464338 209080 464344 209092
rect 445168 209052 464344 209080
rect 445168 209040 445174 209052
rect 464338 209040 464344 209052
rect 464396 209040 464402 209092
rect 372890 208360 372896 208412
rect 372948 208400 372954 208412
rect 373350 208400 373356 208412
rect 372948 208372 373356 208400
rect 372948 208360 372954 208372
rect 373350 208360 373356 208372
rect 373408 208360 373414 208412
rect 445110 208292 445116 208344
rect 445168 208332 445174 208344
rect 449250 208332 449256 208344
rect 445168 208304 449256 208332
rect 445168 208292 445174 208304
rect 449250 208292 449256 208304
rect 449308 208292 449314 208344
rect 370958 208088 370964 208140
rect 371016 208128 371022 208140
rect 373994 208128 374000 208140
rect 371016 208100 374000 208128
rect 371016 208088 371022 208100
rect 373994 208088 374000 208100
rect 374052 208088 374058 208140
rect 445662 207612 445668 207664
rect 445720 207652 445726 207664
rect 454678 207652 454684 207664
rect 445720 207624 454684 207652
rect 445720 207612 445726 207624
rect 454678 207612 454684 207624
rect 454736 207612 454742 207664
rect 181622 207000 181628 207052
rect 181680 207040 181686 207052
rect 197354 207040 197360 207052
rect 181680 207012 197360 207040
rect 181680 207000 181686 207012
rect 197354 207000 197360 207012
rect 197412 207000 197418 207052
rect 516134 206864 516140 206916
rect 516192 206904 516198 206916
rect 528646 206904 528652 206916
rect 516192 206876 528652 206904
rect 516192 206864 516198 206876
rect 528646 206864 528652 206876
rect 528704 206864 528710 206916
rect 515398 206796 515404 206848
rect 515456 206836 515462 206848
rect 580166 206836 580172 206848
rect 515456 206808 580172 206836
rect 515456 206796 515462 206808
rect 580166 206796 580172 206808
rect 580224 206796 580230 206848
rect 302234 206116 302240 206168
rect 302292 206156 302298 206168
rect 304258 206156 304264 206168
rect 302292 206128 304264 206156
rect 302292 206116 302298 206128
rect 304258 206116 304264 206128
rect 304316 206116 304322 206168
rect 444374 205844 444380 205896
rect 444432 205884 444438 205896
rect 448146 205884 448152 205896
rect 444432 205856 448152 205884
rect 444432 205844 444438 205856
rect 448146 205844 448152 205856
rect 448204 205844 448210 205896
rect 516134 205844 516140 205896
rect 516192 205884 516198 205896
rect 517790 205884 517796 205896
rect 516192 205856 517796 205884
rect 516192 205844 516198 205856
rect 517790 205844 517796 205856
rect 517848 205844 517854 205896
rect 444282 205708 444288 205760
rect 444340 205748 444346 205760
rect 444650 205748 444656 205760
rect 444340 205720 444656 205748
rect 444340 205708 444346 205720
rect 444650 205708 444656 205720
rect 444708 205708 444714 205760
rect 180242 205640 180248 205692
rect 180300 205680 180306 205692
rect 197354 205680 197360 205692
rect 180300 205652 197360 205680
rect 180300 205640 180306 205652
rect 197354 205640 197360 205652
rect 197412 205640 197418 205692
rect 443638 205572 443644 205624
rect 443696 205612 443702 205624
rect 444190 205612 444196 205624
rect 443696 205584 444196 205612
rect 443696 205572 443702 205584
rect 444190 205572 444196 205584
rect 444248 205612 444254 205624
rect 447962 205612 447968 205624
rect 444248 205584 447968 205612
rect 444248 205572 444254 205584
rect 447962 205572 447968 205584
rect 448020 205572 448026 205624
rect 442902 205300 442908 205352
rect 442960 205340 442966 205352
rect 446674 205340 446680 205352
rect 442960 205312 446680 205340
rect 442960 205300 442966 205312
rect 446674 205300 446680 205312
rect 446732 205300 446738 205352
rect 516134 204892 516140 204944
rect 516192 204932 516198 204944
rect 516318 204932 516324 204944
rect 516192 204904 516324 204932
rect 516192 204892 516198 204904
rect 516318 204892 516324 204904
rect 516376 204932 516382 204944
rect 525886 204932 525892 204944
rect 516376 204904 525892 204932
rect 516376 204892 516382 204904
rect 525886 204892 525892 204904
rect 525944 204892 525950 204944
rect 444374 204756 444380 204808
rect 444432 204796 444438 204808
rect 447778 204796 447784 204808
rect 444432 204768 447784 204796
rect 444432 204756 444438 204768
rect 447778 204756 447784 204768
rect 447836 204756 447842 204808
rect 516134 204212 516140 204264
rect 516192 204252 516198 204264
rect 524598 204252 524604 204264
rect 516192 204224 524604 204252
rect 516192 204212 516198 204224
rect 524598 204212 524604 204224
rect 524656 204212 524662 204264
rect 442718 203940 442724 203992
rect 442776 203980 442782 203992
rect 446398 203980 446404 203992
rect 442776 203952 446404 203980
rect 442776 203940 442782 203952
rect 446398 203940 446404 203952
rect 446456 203940 446462 203992
rect 442350 203328 442356 203380
rect 442408 203368 442414 203380
rect 446582 203368 446588 203380
rect 442408 203340 446588 203368
rect 442408 203328 442414 203340
rect 446582 203328 446588 203340
rect 446640 203328 446646 203380
rect 173250 202852 173256 202904
rect 173308 202892 173314 202904
rect 198274 202892 198280 202904
rect 173308 202864 198280 202892
rect 173308 202852 173314 202864
rect 198274 202852 198280 202864
rect 198332 202852 198338 202904
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 28258 202824 28264 202836
rect 3476 202796 28264 202824
rect 3476 202784 3482 202796
rect 28258 202784 28264 202796
rect 28316 202784 28322 202836
rect 447226 202784 447232 202836
rect 447284 202824 447290 202836
rect 447870 202824 447876 202836
rect 447284 202796 447876 202824
rect 447284 202784 447290 202796
rect 447870 202784 447876 202796
rect 447928 202784 447934 202836
rect 516134 202784 516140 202836
rect 516192 202824 516198 202836
rect 521746 202824 521752 202836
rect 516192 202796 521752 202824
rect 516192 202784 516198 202796
rect 521746 202784 521752 202796
rect 521804 202784 521810 202836
rect 442902 202716 442908 202768
rect 442960 202756 442966 202768
rect 446490 202756 446496 202768
rect 442960 202728 446496 202756
rect 442960 202716 442966 202728
rect 446490 202716 446496 202728
rect 446548 202716 446554 202768
rect 371602 202308 371608 202360
rect 371660 202348 371666 202360
rect 371878 202348 371884 202360
rect 371660 202320 371884 202348
rect 371660 202308 371666 202320
rect 371878 202308 371884 202320
rect 371936 202308 371942 202360
rect 173158 201492 173164 201544
rect 173216 201532 173222 201544
rect 197354 201532 197360 201544
rect 173216 201504 197360 201532
rect 173216 201492 173222 201504
rect 197354 201492 197360 201504
rect 197412 201492 197418 201544
rect 445662 201492 445668 201544
rect 445720 201532 445726 201544
rect 447226 201532 447232 201544
rect 445720 201504 447232 201532
rect 445720 201492 445726 201504
rect 447226 201492 447232 201504
rect 447284 201492 447290 201544
rect 514662 201220 514668 201272
rect 514720 201260 514726 201272
rect 520642 201260 520648 201272
rect 514720 201232 520648 201260
rect 514720 201220 514726 201232
rect 520642 201220 520648 201232
rect 520700 201220 520706 201272
rect 445202 200064 445208 200116
rect 445260 200104 445266 200116
rect 445386 200104 445392 200116
rect 445260 200076 445392 200104
rect 445260 200064 445266 200076
rect 445386 200064 445392 200076
rect 445444 200064 445450 200116
rect 514202 200064 514208 200116
rect 514260 200104 514266 200116
rect 525794 200104 525800 200116
rect 514260 200076 525800 200104
rect 514260 200064 514266 200076
rect 525794 200064 525800 200076
rect 525852 200064 525858 200116
rect 514110 199996 514116 200048
rect 514168 200036 514174 200048
rect 523034 200036 523040 200048
rect 514168 200008 523040 200036
rect 514168 199996 514174 200008
rect 523034 199996 523040 200008
rect 523092 199996 523098 200048
rect 303430 199384 303436 199436
rect 303488 199424 303494 199436
rect 346302 199424 346308 199436
rect 303488 199396 346308 199424
rect 303488 199384 303494 199396
rect 346302 199384 346308 199396
rect 346360 199384 346366 199436
rect 173434 198704 173440 198756
rect 173492 198744 173498 198756
rect 197538 198744 197544 198756
rect 173492 198716 197544 198744
rect 173492 198704 173498 198716
rect 197538 198704 197544 198716
rect 197596 198704 197602 198756
rect 514110 198636 514116 198688
rect 514168 198676 514174 198688
rect 520274 198676 520280 198688
rect 514168 198648 520280 198676
rect 514168 198636 514174 198648
rect 520274 198636 520280 198648
rect 520332 198636 520338 198688
rect 445294 198024 445300 198076
rect 445352 198064 445358 198076
rect 513558 198064 513564 198076
rect 445352 198036 513564 198064
rect 445352 198024 445358 198036
rect 513558 198024 513564 198036
rect 513616 198024 513622 198076
rect 476482 197956 476488 198008
rect 476540 197996 476546 198008
rect 513374 197996 513380 198008
rect 476540 197968 513380 197996
rect 476540 197956 476546 197968
rect 513374 197956 513380 197968
rect 513432 197956 513438 198008
rect 444926 197752 444932 197804
rect 444984 197792 444990 197804
rect 445294 197792 445300 197804
rect 444984 197764 445300 197792
rect 444984 197752 444990 197764
rect 445294 197752 445300 197764
rect 445352 197752 445358 197804
rect 370958 197616 370964 197668
rect 371016 197656 371022 197668
rect 372614 197656 372620 197668
rect 371016 197628 372620 197656
rect 371016 197616 371022 197628
rect 372614 197616 372620 197628
rect 372672 197656 372678 197668
rect 374086 197656 374092 197668
rect 372672 197628 374092 197656
rect 372672 197616 372678 197628
rect 374086 197616 374092 197628
rect 374144 197616 374150 197668
rect 173342 197344 173348 197396
rect 173400 197384 173406 197396
rect 197354 197384 197360 197396
rect 173400 197356 197360 197384
rect 173400 197344 173406 197356
rect 197354 197344 197360 197356
rect 197412 197344 197418 197396
rect 369118 197344 369124 197396
rect 369176 197384 369182 197396
rect 369302 197384 369308 197396
rect 369176 197356 369308 197384
rect 369176 197344 369182 197356
rect 369302 197344 369308 197356
rect 369360 197344 369366 197396
rect 445294 197344 445300 197396
rect 445352 197384 445358 197396
rect 476482 197384 476488 197396
rect 445352 197356 476488 197384
rect 445352 197344 445358 197356
rect 476482 197344 476488 197356
rect 476540 197384 476546 197396
rect 476758 197384 476764 197396
rect 476540 197356 476764 197384
rect 476540 197344 476546 197356
rect 476758 197344 476764 197356
rect 476816 197344 476822 197396
rect 445754 197276 445760 197328
rect 445812 197316 445818 197328
rect 445812 197288 451274 197316
rect 445812 197276 445818 197288
rect 369854 197208 369860 197260
rect 369912 197248 369918 197260
rect 371142 197248 371148 197260
rect 369912 197220 371148 197248
rect 369912 197208 369918 197220
rect 371142 197208 371148 197220
rect 371200 197248 371206 197260
rect 443362 197248 443368 197260
rect 371200 197220 443368 197248
rect 371200 197208 371206 197220
rect 443362 197208 443368 197220
rect 443420 197208 443426 197260
rect 445386 197208 445392 197260
rect 445444 197248 445450 197260
rect 447134 197248 447140 197260
rect 445444 197220 447140 197248
rect 445444 197208 445450 197220
rect 447134 197208 447140 197220
rect 447192 197208 447198 197260
rect 451246 197248 451274 197288
rect 513282 197276 513288 197328
rect 513340 197316 513346 197328
rect 514938 197316 514944 197328
rect 513340 197288 514944 197316
rect 513340 197276 513346 197288
rect 514938 197276 514944 197288
rect 514996 197276 515002 197328
rect 516502 197248 516508 197260
rect 451246 197220 516508 197248
rect 516502 197208 516508 197220
rect 516560 197208 516566 197260
rect 445202 197140 445208 197192
rect 445260 197180 445266 197192
rect 445478 197180 445484 197192
rect 445260 197152 445484 197180
rect 445260 197140 445266 197152
rect 445478 197140 445484 197152
rect 445536 197180 445542 197192
rect 516318 197180 516324 197192
rect 445536 197152 516324 197180
rect 445536 197140 445542 197152
rect 516318 197140 516324 197152
rect 516376 197140 516382 197192
rect 466914 196800 466920 196852
rect 466972 196840 466978 196852
rect 514202 196840 514208 196852
rect 466972 196812 514208 196840
rect 466972 196800 466978 196812
rect 514202 196800 514208 196812
rect 514260 196800 514266 196852
rect 447134 196664 447140 196716
rect 447192 196704 447198 196716
rect 457438 196704 457444 196716
rect 447192 196676 457444 196704
rect 447192 196664 447198 196676
rect 457438 196664 457444 196676
rect 457496 196704 457502 196716
rect 514110 196704 514116 196716
rect 457496 196676 514116 196704
rect 457496 196664 457502 196676
rect 514110 196664 514116 196676
rect 514168 196664 514174 196716
rect 302786 196596 302792 196648
rect 302844 196636 302850 196648
rect 369854 196636 369860 196648
rect 302844 196608 369860 196636
rect 302844 196596 302850 196608
rect 369854 196596 369860 196608
rect 369912 196596 369918 196648
rect 445570 196596 445576 196648
rect 445628 196636 445634 196648
rect 460198 196636 460204 196648
rect 445628 196608 460204 196636
rect 445628 196596 445634 196608
rect 460198 196596 460204 196608
rect 460256 196636 460262 196648
rect 516134 196636 516140 196648
rect 460256 196608 516140 196636
rect 460256 196596 460262 196608
rect 516134 196596 516140 196608
rect 516192 196596 516198 196648
rect 445754 196052 445760 196104
rect 445812 196092 445818 196104
rect 446490 196092 446496 196104
rect 445812 196064 446496 196092
rect 445812 196052 445818 196064
rect 446490 196052 446496 196064
rect 446548 196052 446554 196104
rect 445662 195984 445668 196036
rect 445720 196024 445726 196036
rect 466914 196024 466920 196036
rect 445720 195996 466920 196024
rect 445720 195984 445726 195996
rect 466914 195984 466920 195996
rect 466972 195984 466978 196036
rect 346302 195304 346308 195356
rect 346360 195344 346366 195356
rect 381538 195344 381544 195356
rect 346360 195316 381544 195344
rect 346360 195304 346366 195316
rect 381538 195304 381544 195316
rect 381596 195344 381602 195356
rect 381596 195316 383654 195344
rect 381596 195304 381602 195316
rect 303338 195236 303344 195288
rect 303396 195276 303402 195288
rect 370314 195276 370320 195288
rect 303396 195248 370320 195276
rect 303396 195236 303402 195248
rect 370314 195236 370320 195248
rect 370372 195236 370378 195288
rect 383626 195276 383654 195316
rect 445938 195276 445944 195288
rect 383626 195248 445944 195276
rect 445938 195236 445944 195248
rect 445996 195236 446002 195288
rect 173526 194556 173532 194608
rect 173584 194596 173590 194608
rect 197538 194596 197544 194608
rect 173584 194568 197544 194596
rect 173584 194556 173590 194568
rect 197538 194556 197544 194568
rect 197596 194556 197602 194608
rect 305638 194488 305644 194540
rect 305696 194528 305702 194540
rect 510890 194528 510896 194540
rect 305696 194500 510896 194528
rect 305696 194488 305702 194500
rect 510890 194488 510896 194500
rect 510948 194488 510954 194540
rect 359458 194420 359464 194472
rect 359516 194460 359522 194472
rect 366910 194460 366916 194472
rect 359516 194432 366916 194460
rect 359516 194420 359522 194432
rect 366910 194420 366916 194432
rect 366968 194420 366974 194472
rect 371970 194420 371976 194472
rect 372028 194460 372034 194472
rect 375374 194460 375380 194472
rect 372028 194432 375380 194460
rect 372028 194420 372034 194432
rect 375374 194420 375380 194432
rect 375432 194460 375438 194472
rect 443270 194460 443276 194472
rect 375432 194432 443276 194460
rect 375432 194420 375438 194432
rect 443270 194420 443276 194432
rect 443328 194420 443334 194472
rect 506842 194420 506848 194472
rect 506900 194460 506906 194472
rect 507762 194460 507768 194472
rect 506900 194432 507768 194460
rect 506900 194420 506906 194432
rect 507762 194420 507768 194432
rect 507820 194460 507826 194472
rect 514754 194460 514760 194472
rect 507820 194432 514760 194460
rect 507820 194420 507826 194432
rect 514754 194420 514760 194432
rect 514812 194420 514818 194472
rect 508866 194352 508872 194404
rect 508924 194392 508930 194404
rect 514846 194392 514852 194404
rect 508924 194364 514852 194392
rect 508924 194352 508930 194364
rect 514846 194352 514852 194364
rect 514904 194352 514910 194404
rect 305730 193808 305736 193860
rect 305788 193848 305794 193860
rect 438946 193848 438952 193860
rect 305788 193820 438952 193848
rect 305788 193808 305794 193820
rect 438946 193808 438952 193820
rect 439004 193808 439010 193860
rect 173618 193196 173624 193248
rect 173676 193236 173682 193248
rect 197354 193236 197360 193248
rect 173676 193208 197360 193236
rect 173676 193196 173682 193208
rect 197354 193196 197360 193208
rect 197412 193196 197418 193248
rect 302602 193196 302608 193248
rect 302660 193236 302666 193248
rect 371050 193236 371056 193248
rect 302660 193208 371056 193236
rect 302660 193196 302666 193208
rect 371050 193196 371056 193208
rect 371108 193236 371114 193248
rect 371970 193236 371976 193248
rect 371108 193208 371976 193236
rect 371108 193196 371114 193208
rect 371970 193196 371976 193208
rect 372028 193196 372034 193248
rect 522298 193128 522304 193180
rect 522356 193168 522362 193180
rect 580166 193168 580172 193180
rect 522356 193140 580172 193168
rect 522356 193128 522362 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 302418 191768 302424 191820
rect 302476 191808 302482 191820
rect 369210 191808 369216 191820
rect 302476 191780 369216 191808
rect 302476 191768 302482 191780
rect 369210 191768 369216 191780
rect 369268 191808 369274 191820
rect 370958 191808 370964 191820
rect 369268 191780 370964 191808
rect 369268 191768 369274 191780
rect 370958 191768 370964 191780
rect 371016 191808 371022 191820
rect 371694 191808 371700 191820
rect 371016 191780 371700 191808
rect 371016 191768 371022 191780
rect 371694 191768 371700 191780
rect 371752 191768 371758 191820
rect 371694 191088 371700 191140
rect 371752 191128 371758 191140
rect 442258 191128 442264 191140
rect 371752 191100 442264 191128
rect 371752 191088 371758 191100
rect 442258 191088 442264 191100
rect 442316 191088 442322 191140
rect 193950 190884 193956 190936
rect 194008 190924 194014 190936
rect 198274 190924 198280 190936
rect 194008 190896 198280 190924
rect 194008 190884 194014 190896
rect 198274 190884 198280 190896
rect 198332 190884 198338 190936
rect 172422 190068 172428 190120
rect 172480 190108 172486 190120
rect 175918 190108 175924 190120
rect 172480 190080 175924 190108
rect 172480 190068 172486 190080
rect 175918 190068 175924 190080
rect 175976 190068 175982 190120
rect 352558 189728 352564 189780
rect 352616 189768 352622 189780
rect 374454 189768 374460 189780
rect 352616 189740 374460 189768
rect 352616 189728 352622 189740
rect 374454 189728 374460 189740
rect 374512 189768 374518 189780
rect 375282 189768 375288 189780
rect 374512 189740 375288 189768
rect 374512 189728 374518 189740
rect 375282 189728 375288 189740
rect 375340 189728 375346 189780
rect 176102 189048 176108 189100
rect 176160 189088 176166 189100
rect 197354 189088 197360 189100
rect 176160 189060 197360 189088
rect 176160 189048 176166 189060
rect 197354 189048 197360 189060
rect 197412 189048 197418 189100
rect 375282 189048 375288 189100
rect 375340 189088 375346 189100
rect 446398 189088 446404 189100
rect 375340 189060 446404 189088
rect 375340 189048 375346 189060
rect 446398 189048 446404 189060
rect 446456 189048 446462 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 155218 189020 155224 189032
rect 3476 188992 155224 189020
rect 3476 188980 3482 188992
rect 155218 188980 155224 188992
rect 155276 188980 155282 189032
rect 172422 188980 172428 189032
rect 172480 189020 172486 189032
rect 181438 189020 181444 189032
rect 172480 188992 181444 189020
rect 172480 188980 172486 188992
rect 181438 188980 181444 188992
rect 181496 188980 181502 189032
rect 172422 187620 172428 187672
rect 172480 187660 172486 187672
rect 188338 187660 188344 187672
rect 172480 187632 188344 187660
rect 172480 187620 172486 187632
rect 188338 187620 188344 187632
rect 188396 187620 188402 187672
rect 376938 187620 376944 187672
rect 376996 187660 377002 187672
rect 443454 187660 443460 187672
rect 376996 187632 443460 187660
rect 376996 187620 377002 187632
rect 443454 187620 443460 187632
rect 443512 187620 443518 187672
rect 303062 186940 303068 186992
rect 303120 186980 303126 186992
rect 303430 186980 303436 186992
rect 303120 186952 303436 186980
rect 303120 186940 303126 186952
rect 303430 186940 303436 186952
rect 303488 186980 303494 186992
rect 376938 186980 376944 186992
rect 303488 186952 376944 186980
rect 303488 186940 303494 186952
rect 376938 186940 376944 186952
rect 376996 186940 377002 186992
rect 174722 186328 174728 186380
rect 174780 186368 174786 186380
rect 197354 186368 197360 186380
rect 174780 186340 197360 186368
rect 174780 186328 174786 186340
rect 197354 186328 197360 186340
rect 197412 186328 197418 186380
rect 172422 186192 172428 186244
rect 172480 186232 172486 186244
rect 180058 186232 180064 186244
rect 172480 186204 180064 186232
rect 172480 186192 172486 186204
rect 180058 186192 180064 186204
rect 180116 186192 180122 186244
rect 196802 184968 196808 185020
rect 196860 185008 196866 185020
rect 198458 185008 198464 185020
rect 196860 184980 198464 185008
rect 196860 184968 196866 184980
rect 198458 184968 198464 184980
rect 198516 184968 198522 185020
rect 172330 184832 172336 184884
rect 172388 184872 172394 184884
rect 193858 184872 193864 184884
rect 172388 184844 193864 184872
rect 172388 184832 172394 184844
rect 193858 184832 193864 184844
rect 193916 184832 193922 184884
rect 302786 184832 302792 184884
rect 302844 184872 302850 184884
rect 376846 184872 376852 184884
rect 302844 184844 376852 184872
rect 302844 184832 302850 184844
rect 376846 184832 376852 184844
rect 376904 184872 376910 184884
rect 378042 184872 378048 184884
rect 376904 184844 378048 184872
rect 376904 184832 376910 184844
rect 378042 184832 378048 184844
rect 378100 184832 378106 184884
rect 172422 184764 172428 184816
rect 172480 184804 172486 184816
rect 186958 184804 186964 184816
rect 172480 184776 186964 184804
rect 172480 184764 172486 184776
rect 186958 184764 186964 184776
rect 187016 184764 187022 184816
rect 378042 184152 378048 184204
rect 378100 184192 378106 184204
rect 399478 184192 399484 184204
rect 378100 184164 399484 184192
rect 378100 184152 378106 184164
rect 399478 184152 399484 184164
rect 399536 184192 399542 184204
rect 442166 184192 442172 184204
rect 399536 184164 442172 184192
rect 399536 184152 399542 184164
rect 442166 184152 442172 184164
rect 442224 184152 442230 184204
rect 172422 183472 172428 183524
rect 172480 183512 172486 183524
rect 184198 183512 184204 183524
rect 172480 183484 184204 183512
rect 172480 183472 172486 183484
rect 184198 183472 184204 183484
rect 184256 183472 184262 183524
rect 178862 182180 178868 182232
rect 178920 182220 178926 182232
rect 197354 182220 197360 182232
rect 178920 182192 197360 182220
rect 178920 182180 178926 182192
rect 197354 182180 197360 182192
rect 197412 182180 197418 182232
rect 172422 182112 172428 182164
rect 172480 182152 172486 182164
rect 182818 182152 182824 182164
rect 172480 182124 182824 182152
rect 172480 182112 172486 182124
rect 182818 182112 182824 182124
rect 182876 182112 182882 182164
rect 302694 182112 302700 182164
rect 302752 182152 302758 182164
rect 377674 182152 377680 182164
rect 302752 182124 377680 182152
rect 302752 182112 302758 182124
rect 377674 182112 377680 182124
rect 377732 182152 377738 182164
rect 378042 182152 378048 182164
rect 377732 182124 378048 182152
rect 377732 182112 377738 182124
rect 378042 182112 378048 182124
rect 378100 182112 378106 182164
rect 378042 181432 378048 181484
rect 378100 181472 378106 181484
rect 395338 181472 395344 181484
rect 378100 181444 395344 181472
rect 378100 181432 378106 181444
rect 395338 181432 395344 181444
rect 395396 181472 395402 181484
rect 443086 181472 443092 181484
rect 395396 181444 443092 181472
rect 395396 181432 395402 181444
rect 443086 181432 443092 181444
rect 443144 181432 443150 181484
rect 195422 180888 195428 180940
rect 195480 180928 195486 180940
rect 198274 180928 198280 180940
rect 195480 180900 198280 180928
rect 195480 180888 195486 180900
rect 198274 180888 198280 180900
rect 198332 180888 198338 180940
rect 172422 180752 172428 180804
rect 172480 180792 172486 180804
rect 181530 180792 181536 180804
rect 172480 180764 181536 180792
rect 172480 180752 172486 180764
rect 181530 180752 181536 180764
rect 181588 180752 181594 180804
rect 373626 179432 373632 179444
rect 304920 179404 373632 179432
rect 304920 179376 304948 179404
rect 373626 179392 373632 179404
rect 373684 179392 373690 179444
rect 303338 179324 303344 179376
rect 303396 179364 303402 179376
rect 304902 179364 304908 179376
rect 303396 179336 304908 179364
rect 303396 179324 303402 179336
rect 304902 179324 304908 179336
rect 304960 179324 304966 179376
rect 536098 179324 536104 179376
rect 536156 179364 536162 179376
rect 580166 179364 580172 179376
rect 536156 179336 580172 179364
rect 536156 179324 536162 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 171134 179188 171140 179240
rect 171192 179228 171198 179240
rect 180150 179228 180156 179240
rect 171192 179200 180156 179228
rect 171192 179188 171198 179200
rect 180150 179188 180156 179200
rect 180208 179188 180214 179240
rect 373534 178644 373540 178696
rect 373592 178684 373598 178696
rect 442258 178684 442264 178696
rect 373592 178656 442264 178684
rect 373592 178644 373598 178656
rect 442258 178644 442264 178656
rect 442316 178644 442322 178696
rect 180334 178032 180340 178084
rect 180392 178072 180398 178084
rect 197354 178072 197360 178084
rect 180392 178044 197360 178072
rect 180392 178032 180398 178044
rect 197354 178032 197360 178044
rect 197412 178032 197418 178084
rect 172238 177964 172244 178016
rect 172296 178004 172302 178016
rect 196618 178004 196624 178016
rect 172296 177976 196624 178004
rect 172296 177964 172302 177976
rect 196618 177964 196624 177976
rect 196676 177964 196682 178016
rect 172422 177896 172428 177948
rect 172480 177936 172486 177948
rect 178770 177936 178776 177948
rect 172480 177908 178776 177936
rect 172480 177896 172486 177908
rect 178770 177896 178776 177908
rect 178828 177896 178834 177948
rect 188338 176672 188344 176724
rect 188396 176712 188402 176724
rect 197354 176712 197360 176724
rect 188396 176684 197360 176712
rect 188396 176672 188402 176684
rect 197354 176672 197360 176684
rect 197412 176672 197418 176724
rect 172238 176604 172244 176656
rect 172296 176644 172302 176656
rect 195238 176644 195244 176656
rect 172296 176616 195244 176644
rect 172296 176604 172302 176616
rect 195238 176604 195244 176616
rect 195296 176604 195302 176656
rect 368382 176604 368388 176656
rect 368440 176644 368446 176656
rect 372798 176644 372804 176656
rect 368440 176616 372804 176644
rect 368440 176604 368446 176616
rect 372798 176604 372804 176616
rect 372856 176644 372862 176656
rect 441982 176644 441988 176656
rect 372856 176616 441988 176644
rect 372856 176604 372862 176616
rect 441982 176604 441988 176616
rect 442040 176604 442046 176656
rect 302234 175244 302240 175296
rect 302292 175284 302298 175296
rect 357250 175284 357256 175296
rect 302292 175256 357256 175284
rect 302292 175244 302298 175256
rect 357250 175244 357256 175256
rect 357308 175284 357314 175296
rect 358078 175284 358084 175296
rect 357308 175256 358084 175284
rect 357308 175244 357314 175256
rect 358078 175244 358084 175256
rect 358136 175244 358142 175296
rect 441982 175244 441988 175296
rect 442040 175284 442046 175296
rect 442350 175284 442356 175296
rect 442040 175256 442356 175284
rect 442040 175244 442046 175256
rect 442350 175244 442356 175256
rect 442408 175244 442414 175296
rect 172422 175176 172428 175228
rect 172480 175216 172486 175228
rect 192570 175216 192576 175228
rect 172480 175188 192576 175216
rect 172480 175176 172486 175188
rect 192570 175176 192576 175188
rect 192628 175176 192634 175228
rect 186958 173884 186964 173936
rect 187016 173924 187022 173936
rect 197722 173924 197728 173936
rect 187016 173896 197728 173924
rect 187016 173884 187022 173896
rect 197722 173884 197728 173896
rect 197780 173884 197786 173936
rect 172422 173816 172428 173868
rect 172480 173856 172486 173868
rect 191190 173856 191196 173868
rect 172480 173828 191196 173856
rect 172480 173816 172486 173828
rect 191190 173816 191196 173828
rect 191248 173816 191254 173868
rect 184198 172524 184204 172576
rect 184256 172564 184262 172576
rect 197354 172564 197360 172576
rect 184256 172536 197360 172564
rect 184256 172524 184262 172536
rect 197354 172524 197360 172536
rect 197412 172524 197418 172576
rect 372430 172524 372436 172576
rect 372488 172564 372494 172576
rect 442718 172564 442724 172576
rect 372488 172536 442724 172564
rect 372488 172524 372494 172536
rect 442718 172524 442724 172536
rect 442776 172564 442782 172576
rect 444742 172564 444748 172576
rect 442776 172536 444748 172564
rect 442776 172524 442782 172536
rect 444742 172524 444748 172536
rect 444800 172524 444806 172576
rect 172422 172388 172428 172440
rect 172480 172428 172486 172440
rect 177390 172428 177396 172440
rect 172480 172400 177396 172428
rect 172480 172388 172486 172400
rect 177390 172388 177396 172400
rect 177448 172388 177454 172440
rect 373442 171776 373448 171828
rect 373500 171816 373506 171828
rect 442442 171816 442448 171828
rect 373500 171788 442448 171816
rect 373500 171776 373506 171788
rect 442442 171776 442448 171788
rect 442500 171776 442506 171828
rect 172422 171028 172428 171080
rect 172480 171068 172486 171080
rect 198090 171068 198096 171080
rect 172480 171040 198096 171068
rect 172480 171028 172486 171040
rect 198090 171028 198096 171040
rect 198148 171028 198154 171080
rect 442626 171028 442632 171080
rect 442684 171068 442690 171080
rect 445110 171068 445116 171080
rect 442684 171040 445116 171068
rect 442684 171028 442690 171040
rect 445110 171028 445116 171040
rect 445168 171028 445174 171080
rect 371234 170484 371240 170536
rect 371292 170524 371298 170536
rect 371878 170524 371884 170536
rect 371292 170496 371884 170524
rect 371292 170484 371298 170496
rect 371878 170484 371884 170496
rect 371936 170484 371942 170536
rect 371234 170348 371240 170400
rect 371292 170388 371298 170400
rect 376018 170388 376024 170400
rect 371292 170360 376024 170388
rect 371292 170348 371298 170360
rect 376018 170348 376024 170360
rect 376076 170388 376082 170400
rect 442626 170388 442632 170400
rect 376076 170360 442632 170388
rect 376076 170348 376082 170360
rect 442626 170348 442632 170360
rect 442684 170348 442690 170400
rect 172238 169668 172244 169720
rect 172296 169708 172302 169720
rect 195330 169708 195336 169720
rect 172296 169680 195336 169708
rect 172296 169668 172302 169680
rect 195330 169668 195336 169680
rect 195388 169668 195394 169720
rect 371694 169260 371700 169312
rect 371752 169300 371758 169312
rect 372430 169300 372436 169312
rect 371752 169272 372436 169300
rect 371752 169260 371758 169272
rect 372430 169260 372436 169272
rect 372488 169260 372494 169312
rect 302786 168988 302792 169040
rect 302844 169028 302850 169040
rect 371694 169028 371700 169040
rect 302844 169000 371700 169028
rect 302844 168988 302850 169000
rect 371694 168988 371700 169000
rect 371752 168988 371758 169040
rect 373718 168308 373724 168360
rect 373776 168348 373782 168360
rect 374362 168348 374368 168360
rect 373776 168320 374368 168348
rect 373776 168308 373782 168320
rect 374362 168308 374368 168320
rect 374420 168348 374426 168360
rect 441798 168348 441804 168360
rect 374420 168320 441804 168348
rect 374420 168308 374426 168320
rect 441798 168308 441804 168320
rect 441856 168348 441862 168360
rect 445110 168348 445116 168360
rect 441856 168320 445116 168348
rect 441856 168308 441862 168320
rect 445110 168308 445116 168320
rect 445168 168308 445174 168360
rect 178770 167628 178776 167680
rect 178828 167668 178834 167680
rect 197446 167668 197452 167680
rect 178828 167640 197452 167668
rect 178828 167628 178834 167640
rect 197446 167628 197452 167640
rect 197504 167628 197510 167680
rect 371878 167628 371884 167680
rect 371936 167668 371942 167680
rect 444834 167668 444840 167680
rect 371936 167640 444840 167668
rect 371936 167628 371942 167640
rect 444834 167628 444840 167640
rect 444892 167628 444898 167680
rect 444834 167288 444840 167340
rect 444892 167328 444898 167340
rect 445018 167328 445024 167340
rect 444892 167300 445024 167328
rect 444892 167288 444898 167300
rect 445018 167288 445024 167300
rect 445076 167288 445082 167340
rect 182818 167016 182824 167068
rect 182876 167056 182882 167068
rect 197354 167056 197360 167068
rect 182876 167028 197360 167056
rect 182876 167016 182882 167028
rect 197354 167016 197360 167028
rect 197412 167016 197418 167068
rect 172422 166948 172428 167000
rect 172480 166988 172486 167000
rect 196710 166988 196716 167000
rect 172480 166960 196716 166988
rect 172480 166948 172486 166960
rect 196710 166948 196716 166960
rect 196768 166948 196774 167000
rect 301498 166948 301504 167000
rect 301556 166988 301562 167000
rect 580166 166988 580172 167000
rect 301556 166960 580172 166988
rect 301556 166948 301562 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 302786 166268 302792 166320
rect 302844 166308 302850 166320
rect 371970 166308 371976 166320
rect 302844 166280 371976 166308
rect 302844 166268 302850 166280
rect 371970 166268 371976 166280
rect 372028 166308 372034 166320
rect 372338 166308 372344 166320
rect 372028 166280 372344 166308
rect 372028 166268 372034 166280
rect 372338 166268 372344 166280
rect 372396 166268 372402 166320
rect 172146 165520 172152 165572
rect 172204 165560 172210 165572
rect 174630 165560 174636 165572
rect 172204 165532 174636 165560
rect 172204 165520 172210 165532
rect 174630 165520 174636 165532
rect 174688 165520 174694 165572
rect 373350 165520 373356 165572
rect 373408 165560 373414 165572
rect 441890 165560 441896 165572
rect 373408 165532 441896 165560
rect 373408 165520 373414 165532
rect 441890 165520 441896 165532
rect 441948 165560 441954 165572
rect 442994 165560 443000 165572
rect 441948 165532 443000 165560
rect 441948 165520 441954 165532
rect 442994 165520 443000 165532
rect 443052 165520 443058 165572
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 11698 164200 11704 164212
rect 3292 164172 11704 164200
rect 3292 164160 3298 164172
rect 11698 164160 11704 164172
rect 11756 164160 11762 164212
rect 172238 164160 172244 164212
rect 172296 164200 172302 164212
rect 198734 164200 198740 164212
rect 172296 164172 198740 164200
rect 172296 164160 172302 164172
rect 198734 164160 198740 164172
rect 198792 164160 198798 164212
rect 369026 164160 369032 164212
rect 369084 164200 369090 164212
rect 371234 164200 371240 164212
rect 369084 164172 371240 164200
rect 369084 164160 369090 164172
rect 371234 164160 371240 164172
rect 371292 164160 371298 164212
rect 444650 163752 444656 163804
rect 444708 163792 444714 163804
rect 445294 163792 445300 163804
rect 444708 163764 445300 163792
rect 444708 163752 444714 163764
rect 445294 163752 445300 163764
rect 445352 163752 445358 163804
rect 171778 163616 171784 163668
rect 171836 163656 171842 163668
rect 180334 163656 180340 163668
rect 171836 163628 180340 163656
rect 171836 163616 171842 163628
rect 180334 163616 180340 163628
rect 180392 163616 180398 163668
rect 371970 163480 371976 163532
rect 372028 163520 372034 163532
rect 372338 163520 372344 163532
rect 372028 163492 372344 163520
rect 372028 163480 372034 163492
rect 372338 163480 372344 163492
rect 372396 163520 372402 163532
rect 444650 163520 444656 163532
rect 372396 163492 444656 163520
rect 372396 163480 372402 163492
rect 444650 163480 444656 163492
rect 444708 163480 444714 163532
rect 180058 162868 180064 162920
rect 180116 162908 180122 162920
rect 197538 162908 197544 162920
rect 180116 162880 197544 162908
rect 180116 162868 180122 162880
rect 197538 162868 197544 162880
rect 197596 162868 197602 162920
rect 302786 162868 302792 162920
rect 302844 162908 302850 162920
rect 369026 162908 369032 162920
rect 302844 162880 369032 162908
rect 302844 162868 302850 162880
rect 369026 162868 369032 162880
rect 369084 162868 369090 162920
rect 442902 162800 442908 162852
rect 442960 162840 442966 162852
rect 445202 162840 445208 162852
rect 442960 162812 445208 162840
rect 442960 162800 442966 162812
rect 445202 162800 445208 162812
rect 445260 162800 445266 162852
rect 181438 162120 181444 162172
rect 181496 162160 181502 162172
rect 198458 162160 198464 162172
rect 181496 162132 198464 162160
rect 181496 162120 181502 162132
rect 198458 162120 198464 162132
rect 198516 162120 198522 162172
rect 372246 161440 372252 161492
rect 372304 161480 372310 161492
rect 442902 161480 442908 161492
rect 372304 161452 442908 161480
rect 372304 161440 372310 161452
rect 442902 161440 442908 161452
rect 442960 161440 442966 161492
rect 172422 161236 172428 161288
rect 172480 161276 172486 161288
rect 176010 161276 176016 161288
rect 172480 161248 176016 161276
rect 172480 161236 172486 161248
rect 176010 161236 176016 161248
rect 176068 161236 176074 161288
rect 445846 160828 445852 160880
rect 445904 160868 445910 160880
rect 446490 160868 446496 160880
rect 445904 160840 446496 160868
rect 445904 160828 445910 160840
rect 446490 160828 446496 160840
rect 446548 160828 446554 160880
rect 169202 160692 169208 160744
rect 169260 160732 169266 160744
rect 178678 160732 178684 160744
rect 169260 160704 178684 160732
rect 169260 160692 169266 160704
rect 178678 160692 178684 160704
rect 178736 160692 178742 160744
rect 373258 160692 373264 160744
rect 373316 160732 373322 160744
rect 445846 160732 445852 160744
rect 373316 160704 445852 160732
rect 373316 160692 373322 160704
rect 445846 160692 445852 160704
rect 445904 160692 445910 160744
rect 177390 158720 177396 158772
rect 177448 158760 177454 158772
rect 197538 158760 197544 158772
rect 177448 158732 197544 158760
rect 177448 158720 177454 158732
rect 197538 158720 197544 158732
rect 197596 158720 197602 158772
rect 302510 158720 302516 158772
rect 302568 158760 302574 158772
rect 302568 158732 371280 158760
rect 302568 158720 302574 158732
rect 166902 158652 166908 158704
rect 166960 158692 166966 158704
rect 170398 158692 170404 158704
rect 166960 158664 170404 158692
rect 166960 158652 166966 158664
rect 170398 158652 170404 158664
rect 170456 158652 170462 158704
rect 371252 158692 371280 158732
rect 374178 158692 374184 158704
rect 371252 158664 374184 158692
rect 374178 158652 374184 158664
rect 374236 158652 374242 158704
rect 164878 158584 164884 158636
rect 164936 158624 164942 158636
rect 170490 158624 170496 158636
rect 164936 158596 170496 158624
rect 164936 158584 164942 158596
rect 170490 158584 170496 158596
rect 170548 158584 170554 158636
rect 162854 158516 162860 158568
rect 162912 158556 162918 158568
rect 174538 158556 174544 158568
rect 162912 158528 174544 158556
rect 162912 158516 162918 158528
rect 174538 158516 174544 158528
rect 174596 158516 174602 158568
rect 302878 157972 302884 158024
rect 302936 158012 302942 158024
rect 369394 158012 369400 158024
rect 302936 157984 369400 158012
rect 302936 157972 302942 157984
rect 369394 157972 369400 157984
rect 369452 157972 369458 158024
rect 374178 157972 374184 158024
rect 374236 158012 374242 158024
rect 443086 158012 443092 158024
rect 374236 157984 443092 158012
rect 374236 157972 374242 157984
rect 443086 157972 443092 157984
rect 443144 158012 443150 158024
rect 443638 158012 443644 158024
rect 443144 157984 443644 158012
rect 443144 157972 443150 157984
rect 443638 157972 443644 157984
rect 443696 157972 443702 158024
rect 175918 157360 175924 157412
rect 175976 157400 175982 157412
rect 197354 157400 197360 157412
rect 175976 157372 197360 157400
rect 175976 157360 175982 157372
rect 197354 157360 197360 157372
rect 197412 157360 197418 157412
rect 171962 156612 171968 156664
rect 172020 156652 172026 156664
rect 188338 156652 188344 156664
rect 172020 156624 188344 156652
rect 172020 156612 172026 156624
rect 188338 156612 188344 156624
rect 188396 156612 188402 156664
rect 369854 156612 369860 156664
rect 369912 156652 369918 156664
rect 374270 156652 374276 156664
rect 369912 156624 374276 156652
rect 369912 156612 369918 156624
rect 374270 156612 374276 156624
rect 374328 156652 374334 156664
rect 445202 156652 445208 156664
rect 374328 156624 445208 156652
rect 374328 156612 374334 156624
rect 445202 156612 445208 156624
rect 445260 156612 445266 156664
rect 393958 156476 393964 156528
rect 394016 156516 394022 156528
rect 394602 156516 394608 156528
rect 394016 156488 394608 156516
rect 394016 156476 394022 156488
rect 394602 156476 394608 156488
rect 394660 156476 394666 156528
rect 394602 156204 394608 156256
rect 394660 156244 394666 156256
rect 513374 156244 513380 156256
rect 394660 156216 513380 156244
rect 394660 156204 394666 156216
rect 513374 156204 513380 156216
rect 513432 156204 513438 156256
rect 370498 156136 370504 156188
rect 370556 156176 370562 156188
rect 371050 156176 371056 156188
rect 370556 156148 371056 156176
rect 370556 156136 370562 156148
rect 371050 156136 371056 156148
rect 371108 156176 371114 156188
rect 515030 156176 515036 156188
rect 371108 156148 515036 156176
rect 371108 156136 371114 156148
rect 515030 156136 515036 156148
rect 515088 156136 515094 156188
rect 370590 156068 370596 156120
rect 370648 156108 370654 156120
rect 371142 156108 371148 156120
rect 370648 156080 371148 156108
rect 370648 156068 370654 156080
rect 371142 156068 371148 156080
rect 371200 156108 371206 156120
rect 515122 156108 515128 156120
rect 371200 156080 515128 156108
rect 371200 156068 371206 156080
rect 515122 156068 515128 156080
rect 515180 156068 515186 156120
rect 370130 156000 370136 156052
rect 370188 156040 370194 156052
rect 370958 156040 370964 156052
rect 370188 156012 370964 156040
rect 370188 156000 370194 156012
rect 370958 156000 370964 156012
rect 371016 156040 371022 156052
rect 515306 156040 515312 156052
rect 371016 156012 515312 156040
rect 371016 156000 371022 156012
rect 515306 156000 515312 156012
rect 515364 156000 515370 156052
rect 369394 155932 369400 155984
rect 369452 155972 369458 155984
rect 516962 155972 516968 155984
rect 369452 155944 516968 155972
rect 369452 155932 369458 155944
rect 516962 155932 516968 155944
rect 517020 155932 517026 155984
rect 441614 155360 441620 155372
rect 431926 155332 441620 155360
rect 302970 155184 302976 155236
rect 303028 155224 303034 155236
rect 370222 155224 370228 155236
rect 303028 155196 370228 155224
rect 303028 155184 303034 155196
rect 370222 155184 370228 155196
rect 370280 155184 370286 155236
rect 374638 155184 374644 155236
rect 374696 155224 374702 155236
rect 431926 155224 431954 155332
rect 441614 155320 441620 155332
rect 441672 155320 441678 155372
rect 507762 155252 507768 155304
rect 507820 155292 507826 155304
rect 514018 155292 514024 155304
rect 507820 155264 514024 155292
rect 507820 155252 507826 155264
rect 514018 155252 514024 155264
rect 514076 155252 514082 155304
rect 374696 155196 431954 155224
rect 374696 155184 374702 155196
rect 468478 155184 468484 155236
rect 468536 155224 468542 155236
rect 516594 155224 516600 155236
rect 468536 155196 516600 155224
rect 468536 155184 468542 155196
rect 516594 155184 516600 155196
rect 516652 155184 516658 155236
rect 370222 154640 370228 154692
rect 370280 154680 370286 154692
rect 370280 154652 373994 154680
rect 370280 154640 370286 154652
rect 174538 154572 174544 154624
rect 174596 154612 174602 154624
rect 197538 154612 197544 154624
rect 174596 154584 197544 154612
rect 174596 154572 174602 154584
rect 197538 154572 197544 154584
rect 197596 154572 197602 154624
rect 373966 154612 373994 154652
rect 515214 154612 515220 154624
rect 373966 154584 515220 154612
rect 515214 154572 515220 154584
rect 515272 154572 515278 154624
rect 172330 154504 172336 154556
rect 172388 154544 172394 154556
rect 188430 154544 188436 154556
rect 172388 154516 188436 154544
rect 172388 154504 172394 154516
rect 188430 154504 188436 154516
rect 188488 154504 188494 154556
rect 368382 154504 368388 154556
rect 368440 154544 368446 154556
rect 369670 154544 369676 154556
rect 368440 154516 369676 154544
rect 368440 154504 368446 154516
rect 369670 154504 369676 154516
rect 369728 154504 369734 154556
rect 373626 154504 373632 154556
rect 373684 154544 373690 154556
rect 441798 154544 441804 154556
rect 373684 154516 441804 154544
rect 373684 154504 373690 154516
rect 441798 154504 441804 154516
rect 441856 154544 441862 154556
rect 444558 154544 444564 154556
rect 441856 154516 444564 154544
rect 441856 154504 441862 154516
rect 444558 154504 444564 154516
rect 444616 154544 444622 154556
rect 444742 154544 444748 154556
rect 444616 154516 444748 154544
rect 444616 154504 444622 154516
rect 444742 154504 444748 154516
rect 444800 154504 444806 154556
rect 445202 154504 445208 154556
rect 445260 154544 445266 154556
rect 459738 154544 459744 154556
rect 445260 154516 459744 154544
rect 445260 154504 445266 154516
rect 459738 154504 459744 154516
rect 459796 154544 459802 154556
rect 460198 154544 460204 154556
rect 459796 154516 460204 154544
rect 459796 154504 459802 154516
rect 460198 154504 460204 154516
rect 460256 154504 460262 154556
rect 172238 154436 172244 154488
rect 172296 154476 172302 154488
rect 187050 154476 187056 154488
rect 172296 154448 187056 154476
rect 172296 154436 172302 154448
rect 187050 154436 187056 154448
rect 187108 154436 187114 154488
rect 442442 154436 442448 154488
rect 442500 154476 442506 154488
rect 445570 154476 445576 154488
rect 442500 154448 445576 154476
rect 442500 154436 442506 154448
rect 445570 154436 445576 154448
rect 445628 154436 445634 154488
rect 442350 154368 442356 154420
rect 442408 154408 442414 154420
rect 444650 154408 444656 154420
rect 442408 154380 444656 154408
rect 442408 154368 442414 154380
rect 444650 154368 444656 154380
rect 444708 154368 444714 154420
rect 441614 154300 441620 154352
rect 441672 154340 441678 154352
rect 444834 154340 444840 154352
rect 441672 154312 444840 154340
rect 441672 154300 441678 154312
rect 444834 154300 444840 154312
rect 444892 154300 444898 154352
rect 437382 154164 437388 154216
rect 437440 154204 437446 154216
rect 441706 154204 441712 154216
rect 437440 154176 441712 154204
rect 437440 154164 437446 154176
rect 441706 154164 441712 154176
rect 441764 154164 441770 154216
rect 489178 154164 489184 154216
rect 489236 154204 489242 154216
rect 514110 154204 514116 154216
rect 489236 154176 514116 154204
rect 489236 154164 489242 154176
rect 514110 154164 514116 154176
rect 514168 154164 514174 154216
rect 485038 154096 485044 154148
rect 485096 154136 485102 154148
rect 513650 154136 513656 154148
rect 485096 154108 513656 154136
rect 485096 154096 485102 154108
rect 513650 154096 513656 154108
rect 513708 154096 513714 154148
rect 482278 154028 482284 154080
rect 482336 154068 482342 154080
rect 513742 154068 513748 154080
rect 482336 154040 513748 154068
rect 482336 154028 482342 154040
rect 513742 154028 513748 154040
rect 513800 154028 513806 154080
rect 359642 153960 359648 154012
rect 359700 154000 359706 154012
rect 368382 154000 368388 154012
rect 359700 153972 368388 154000
rect 359700 153960 359706 153972
rect 368382 153960 368388 153972
rect 368440 153960 368446 154012
rect 459738 153960 459744 154012
rect 459796 154000 459802 154012
rect 513190 154000 513196 154012
rect 459796 153972 513196 154000
rect 459796 153960 459802 153972
rect 513190 153960 513196 153972
rect 513248 153960 513254 154012
rect 302786 153892 302792 153944
rect 302844 153932 302850 153944
rect 370038 153932 370044 153944
rect 302844 153904 370044 153932
rect 302844 153892 302850 153904
rect 370038 153892 370044 153904
rect 370096 153892 370102 153944
rect 446398 153892 446404 153944
rect 446456 153932 446462 153944
rect 516778 153932 516784 153944
rect 446456 153904 516784 153932
rect 446456 153892 446462 153904
rect 516778 153892 516784 153904
rect 516836 153892 516842 153944
rect 303522 153824 303528 153876
rect 303580 153864 303586 153876
rect 372614 153864 372620 153876
rect 303580 153836 372620 153864
rect 303580 153824 303586 153836
rect 372614 153824 372620 153836
rect 372672 153824 372678 153876
rect 431862 153824 431868 153876
rect 431920 153864 431926 153876
rect 434714 153864 434720 153876
rect 431920 153836 434720 153864
rect 431920 153824 431926 153836
rect 434714 153824 434720 153836
rect 434772 153824 434778 153876
rect 444742 153824 444748 153876
rect 444800 153864 444806 153876
rect 515398 153864 515404 153876
rect 444800 153836 515404 153864
rect 444800 153824 444806 153836
rect 515398 153824 515404 153836
rect 515456 153824 515462 153876
rect 445294 153756 445300 153808
rect 445352 153796 445358 153808
rect 514386 153796 514392 153808
rect 445352 153768 514392 153796
rect 445352 153756 445358 153768
rect 514386 153756 514392 153768
rect 514444 153756 514450 153808
rect 445110 153688 445116 153740
rect 445168 153728 445174 153740
rect 514570 153728 514576 153740
rect 445168 153700 514576 153728
rect 445168 153688 445174 153700
rect 514570 153688 514576 153700
rect 514628 153688 514634 153740
rect 444650 153620 444656 153672
rect 444708 153660 444714 153672
rect 513834 153660 513840 153672
rect 444708 153632 513840 153660
rect 444708 153620 444714 153632
rect 513834 153620 513840 153632
rect 513892 153620 513898 153672
rect 444834 153552 444840 153604
rect 444892 153592 444898 153604
rect 514478 153592 514484 153604
rect 444892 153564 514484 153592
rect 444892 153552 444898 153564
rect 514478 153552 514484 153564
rect 514536 153552 514542 153604
rect 442258 153484 442264 153536
rect 442316 153524 442322 153536
rect 514202 153524 514208 153536
rect 442316 153496 514208 153524
rect 442316 153484 442322 153496
rect 514202 153484 514208 153496
rect 514260 153484 514266 153536
rect 445570 153416 445576 153468
rect 445628 153456 445634 153468
rect 514294 153456 514300 153468
rect 445628 153428 514300 153456
rect 445628 153416 445634 153428
rect 514294 153416 514300 153428
rect 514352 153416 514358 153468
rect 443086 153348 443092 153400
rect 443144 153388 443150 153400
rect 514754 153388 514760 153400
rect 443144 153360 514760 153388
rect 443144 153348 443150 153360
rect 514754 153348 514760 153360
rect 514812 153348 514818 153400
rect 358998 153280 359004 153332
rect 359056 153320 359062 153332
rect 359056 153292 372568 153320
rect 359056 153280 359062 153292
rect 188338 153212 188344 153264
rect 188396 153252 188402 153264
rect 197354 153252 197360 153264
rect 188396 153224 197360 153252
rect 188396 153212 188402 153224
rect 197354 153212 197360 153224
rect 197412 153212 197418 153264
rect 302694 153212 302700 153264
rect 302752 153252 302758 153264
rect 369854 153252 369860 153264
rect 302752 153224 369860 153252
rect 302752 153212 302758 153224
rect 369854 153212 369860 153224
rect 369912 153212 369918 153264
rect 172422 153144 172428 153196
rect 172480 153184 172486 153196
rect 184290 153184 184296 153196
rect 172480 153156 184296 153184
rect 172480 153144 172486 153156
rect 184290 153144 184296 153156
rect 184348 153144 184354 153196
rect 369210 153144 369216 153196
rect 369268 153184 369274 153196
rect 372430 153184 372436 153196
rect 369268 153156 372436 153184
rect 369268 153144 369274 153156
rect 372430 153144 372436 153156
rect 372488 153144 372494 153196
rect 372540 153184 372568 153292
rect 431310 153280 431316 153332
rect 431368 153320 431374 153332
rect 514662 153320 514668 153332
rect 431368 153292 514668 153320
rect 431368 153280 431374 153292
rect 514662 153280 514668 153292
rect 514720 153280 514726 153332
rect 372614 153212 372620 153264
rect 372672 153252 372678 153264
rect 372982 153252 372988 153264
rect 372672 153224 372988 153252
rect 372672 153212 372678 153224
rect 372982 153212 372988 153224
rect 373040 153252 373046 153264
rect 515582 153252 515588 153264
rect 373040 153224 515588 153252
rect 373040 153212 373046 153224
rect 515582 153212 515588 153224
rect 515640 153212 515646 153264
rect 373718 153184 373724 153196
rect 372540 153156 373724 153184
rect 373718 153144 373724 153156
rect 373776 153144 373782 153196
rect 479518 153144 479524 153196
rect 479576 153184 479582 153196
rect 513282 153184 513288 153196
rect 479576 153156 513288 153184
rect 479576 153144 479582 153156
rect 513282 153144 513288 153156
rect 513340 153144 513346 153196
rect 520918 153144 520924 153196
rect 520976 153184 520982 153196
rect 580166 153184 580172 153196
rect 520976 153156 580172 153184
rect 520976 153144 520982 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 172330 153076 172336 153128
rect 172388 153116 172394 153128
rect 182910 153116 182916 153128
rect 172388 153088 182916 153116
rect 172388 153076 172394 153088
rect 182910 153076 182916 153088
rect 182968 153076 182974 153128
rect 370038 153076 370044 153128
rect 370096 153116 370102 153128
rect 372614 153116 372620 153128
rect 370096 153088 372620 153116
rect 370096 153076 370102 153088
rect 372614 153076 372620 153088
rect 372672 153116 372678 153128
rect 373534 153116 373540 153128
rect 372672 153088 373540 153116
rect 372672 153076 372678 153088
rect 373534 153076 373540 153088
rect 373592 153076 373598 153128
rect 493318 153076 493324 153128
rect 493376 153116 493382 153128
rect 513466 153116 513472 153128
rect 493376 153088 513472 153116
rect 493376 153076 493382 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 516226 153076 516232 153128
rect 516284 153116 516290 153128
rect 528830 153116 528836 153128
rect 516284 153088 528836 153116
rect 516284 153076 516290 153088
rect 528830 153076 528836 153088
rect 528888 153076 528894 153128
rect 342162 153008 342168 153060
rect 342220 153048 342226 153060
rect 371234 153048 371240 153060
rect 342220 153020 371240 153048
rect 342220 153008 342226 153020
rect 371234 153008 371240 153020
rect 371292 153008 371298 153060
rect 516134 153008 516140 153060
rect 516192 153048 516198 153060
rect 518894 153048 518900 153060
rect 516192 153020 518900 153048
rect 516192 153008 516198 153020
rect 518894 153008 518900 153020
rect 518952 153008 518958 153060
rect 357342 152940 357348 152992
rect 357400 152980 357406 152992
rect 369486 152980 369492 152992
rect 357400 152952 369492 152980
rect 357400 152940 357406 152952
rect 369486 152940 369492 152952
rect 369544 152940 369550 152992
rect 307662 152872 307668 152924
rect 307720 152912 307726 152924
rect 369578 152912 369584 152924
rect 307720 152884 369584 152912
rect 307720 152872 307726 152884
rect 369578 152872 369584 152884
rect 369636 152872 369642 152924
rect 497458 152872 497464 152924
rect 497516 152912 497522 152924
rect 516686 152912 516692 152924
rect 497516 152884 516692 152912
rect 497516 152872 497522 152884
rect 516686 152872 516692 152884
rect 516744 152872 516750 152924
rect 313182 152804 313188 152856
rect 313240 152844 313246 152856
rect 369302 152844 369308 152856
rect 313240 152816 369308 152844
rect 313240 152804 313246 152816
rect 369302 152804 369308 152816
rect 369360 152804 369366 152856
rect 494698 152804 494704 152856
rect 494756 152844 494762 152856
rect 516502 152844 516508 152856
rect 494756 152816 516508 152844
rect 494756 152804 494762 152816
rect 516502 152804 516508 152816
rect 516560 152804 516566 152856
rect 357250 152736 357256 152788
rect 357308 152776 357314 152788
rect 372706 152776 372712 152788
rect 357308 152748 372712 152776
rect 357308 152736 357314 152748
rect 372706 152736 372712 152748
rect 372764 152736 372770 152788
rect 490558 152736 490564 152788
rect 490616 152776 490622 152788
rect 513374 152776 513380 152788
rect 490616 152748 513380 152776
rect 490616 152736 490622 152748
rect 513374 152736 513380 152748
rect 513432 152736 513438 152788
rect 340782 152668 340788 152720
rect 340840 152708 340846 152720
rect 371234 152708 371240 152720
rect 340840 152680 371240 152708
rect 340840 152668 340846 152680
rect 371234 152668 371240 152680
rect 371292 152668 371298 152720
rect 475378 152668 475384 152720
rect 475436 152708 475442 152720
rect 516318 152708 516324 152720
rect 475436 152680 516324 152708
rect 475436 152668 475442 152680
rect 516318 152668 516324 152680
rect 516376 152668 516382 152720
rect 303062 152600 303068 152652
rect 303120 152640 303126 152652
rect 369210 152640 369216 152652
rect 303120 152612 369216 152640
rect 303120 152600 303126 152612
rect 369210 152600 369216 152612
rect 369268 152600 369274 152652
rect 472618 152600 472624 152652
rect 472676 152640 472682 152652
rect 472676 152612 516180 152640
rect 472676 152600 472682 152612
rect 516152 152584 516180 152612
rect 302786 152532 302792 152584
rect 302844 152572 302850 152584
rect 370038 152572 370044 152584
rect 302844 152544 370044 152572
rect 302844 152532 302850 152544
rect 370038 152532 370044 152544
rect 370096 152572 370102 152584
rect 374638 152572 374644 152584
rect 370096 152544 374644 152572
rect 370096 152532 370102 152544
rect 374638 152532 374644 152544
rect 374696 152532 374702 152584
rect 471238 152532 471244 152584
rect 471296 152572 471302 152584
rect 471296 152544 514064 152572
rect 471296 152532 471302 152544
rect 303430 152464 303436 152516
rect 303488 152504 303494 152516
rect 372890 152504 372896 152516
rect 303488 152476 372896 152504
rect 303488 152464 303494 152476
rect 372890 152464 372896 152476
rect 372948 152464 372954 152516
rect 445662 152464 445668 152516
rect 445720 152504 445726 152516
rect 450538 152504 450544 152516
rect 445720 152476 450544 152504
rect 445720 152464 445726 152476
rect 450538 152464 450544 152476
rect 450596 152504 450602 152516
rect 514036 152504 514064 152544
rect 516134 152532 516140 152584
rect 516192 152532 516198 152584
rect 516410 152504 516416 152516
rect 450596 152476 509234 152504
rect 514036 152476 516416 152504
rect 450596 152464 450602 152476
rect 509206 152164 509234 152476
rect 516410 152464 516416 152476
rect 516468 152464 516474 152516
rect 513926 152164 513932 152176
rect 509206 152136 513932 152164
rect 513926 152124 513932 152136
rect 513984 152124 513990 152176
rect 442718 152056 442724 152108
rect 442776 152096 442782 152108
rect 514938 152096 514944 152108
rect 442776 152068 514944 152096
rect 442776 152056 442782 152068
rect 514938 152056 514944 152068
rect 514996 152056 515002 152108
rect 372706 151988 372712 152040
rect 372764 152028 372770 152040
rect 441798 152028 441804 152040
rect 372764 152000 441804 152028
rect 372764 151988 372770 152000
rect 441798 151988 441804 152000
rect 441856 151988 441862 152040
rect 444742 151988 444748 152040
rect 444800 152028 444806 152040
rect 514846 152028 514852 152040
rect 444800 152000 514852 152028
rect 444800 151988 444806 152000
rect 514846 151988 514852 152000
rect 514904 151988 514910 152040
rect 431402 151920 431408 151972
rect 431460 151960 431466 151972
rect 513098 151960 513104 151972
rect 431460 151932 513104 151960
rect 431460 151920 431466 151932
rect 513098 151920 513104 151932
rect 513156 151920 513162 151972
rect 516502 151920 516508 151972
rect 516560 151920 516566 151972
rect 359550 151852 359556 151904
rect 359608 151892 359614 151904
rect 359608 151864 369808 151892
rect 359608 151852 359614 151864
rect 369780 151768 369808 151864
rect 372890 151852 372896 151904
rect 372948 151892 372954 151904
rect 515490 151892 515496 151904
rect 372948 151864 515496 151892
rect 372948 151852 372954 151864
rect 515490 151852 515496 151864
rect 515548 151852 515554 151904
rect 516318 151852 516324 151904
rect 516376 151892 516382 151904
rect 516520 151892 516548 151920
rect 516376 151864 516548 151892
rect 516376 151852 516382 151864
rect 442626 151784 442632 151836
rect 442684 151824 442690 151836
rect 444190 151824 444196 151836
rect 442684 151796 444196 151824
rect 442684 151784 442690 151796
rect 444190 151784 444196 151796
rect 444248 151784 444254 151836
rect 516502 151784 516508 151836
rect 516560 151824 516566 151836
rect 516962 151824 516968 151836
rect 516560 151796 516968 151824
rect 516560 151784 516566 151796
rect 516962 151784 516968 151796
rect 517020 151784 517026 151836
rect 171686 151716 171692 151768
rect 171744 151756 171750 151768
rect 181622 151756 181628 151768
rect 171744 151728 181628 151756
rect 171744 151716 171750 151728
rect 181622 151716 181628 151728
rect 181680 151716 181686 151768
rect 302786 151716 302792 151768
rect 302844 151756 302850 151768
rect 358998 151756 359004 151768
rect 302844 151728 359004 151756
rect 302844 151716 302850 151728
rect 358998 151716 359004 151728
rect 359056 151716 359062 151768
rect 369762 151716 369768 151768
rect 369820 151756 369826 151768
rect 373442 151756 373448 151768
rect 369820 151728 373448 151756
rect 369820 151716 369826 151728
rect 373442 151716 373448 151728
rect 373500 151716 373506 151768
rect 514110 151716 514116 151768
rect 514168 151756 514174 151768
rect 514168 151728 514340 151756
rect 514168 151716 514174 151728
rect 444374 151648 444380 151700
rect 444432 151688 444438 151700
rect 444742 151688 444748 151700
rect 444432 151660 444748 151688
rect 444432 151648 444438 151660
rect 444742 151648 444748 151660
rect 444800 151648 444806 151700
rect 514202 151648 514208 151700
rect 514260 151648 514266 151700
rect 513558 151580 513564 151632
rect 513616 151620 513622 151632
rect 514220 151620 514248 151648
rect 513616 151592 514248 151620
rect 513616 151580 513622 151592
rect 514312 151496 514340 151728
rect 514386 151648 514392 151700
rect 514444 151648 514450 151700
rect 171502 151444 171508 151496
rect 171560 151484 171566 151496
rect 180242 151484 180248 151496
rect 171560 151456 180248 151484
rect 171560 151444 171566 151456
rect 180242 151444 180248 151456
rect 180300 151444 180306 151496
rect 514294 151444 514300 151496
rect 514352 151444 514358 151496
rect 514294 150628 514300 150680
rect 514352 150668 514358 150680
rect 514404 150668 514432 151648
rect 514352 150640 514432 150668
rect 514352 150628 514358 150640
rect 171594 150560 171600 150612
rect 171652 150600 171658 150612
rect 173250 150600 173256 150612
rect 171652 150572 173256 150600
rect 171652 150560 171658 150572
rect 173250 150560 173256 150572
rect 173308 150560 173314 150612
rect 187050 150424 187056 150476
rect 187108 150464 187114 150476
rect 197538 150464 197544 150476
rect 187108 150436 197544 150464
rect 187108 150424 187114 150436
rect 197538 150424 197544 150436
rect 197596 150424 197602 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 29638 150396 29644 150408
rect 3476 150368 29644 150396
rect 3476 150356 3482 150368
rect 29638 150356 29644 150368
rect 29696 150356 29702 150408
rect 171686 150356 171692 150408
rect 171744 150396 171750 150408
rect 173158 150396 173164 150408
rect 171744 150368 173164 150396
rect 171744 150356 171750 150368
rect 173158 150356 173164 150368
rect 173216 150356 173222 150408
rect 171686 149404 171692 149456
rect 171744 149444 171750 149456
rect 173434 149444 173440 149456
rect 171744 149416 173440 149444
rect 171744 149404 171750 149416
rect 173434 149404 173440 149416
rect 173492 149404 173498 149456
rect 184290 149064 184296 149116
rect 184348 149104 184354 149116
rect 197354 149104 197360 149116
rect 184348 149076 197360 149104
rect 184348 149064 184354 149076
rect 197354 149064 197360 149076
rect 197412 149064 197418 149116
rect 172238 148860 172244 148912
rect 172296 148900 172302 148912
rect 173342 148900 173348 148912
rect 172296 148872 173348 148900
rect 172296 148860 172302 148872
rect 173342 148860 173348 148872
rect 173400 148860 173406 148912
rect 171686 148792 171692 148844
rect 171744 148832 171750 148844
rect 173526 148832 173532 148844
rect 171744 148804 173532 148832
rect 171744 148792 171750 148804
rect 173526 148792 173532 148804
rect 173584 148792 173590 148844
rect 173158 148316 173164 148368
rect 173216 148356 173222 148368
rect 198090 148356 198096 148368
rect 173216 148328 198096 148356
rect 173216 148316 173222 148328
rect 198090 148316 198096 148328
rect 198148 148316 198154 148368
rect 371326 148248 371332 148300
rect 371384 148288 371390 148300
rect 375466 148288 375472 148300
rect 371384 148260 375472 148288
rect 371384 148248 371390 148260
rect 375466 148248 375472 148260
rect 375524 148248 375530 148300
rect 171502 147840 171508 147892
rect 171560 147880 171566 147892
rect 173618 147880 173624 147892
rect 171560 147852 173624 147880
rect 171560 147840 171566 147852
rect 173618 147840 173624 147852
rect 173676 147840 173682 147892
rect 172422 147568 172428 147620
rect 172480 147608 172486 147620
rect 193950 147608 193956 147620
rect 172480 147580 193956 147608
rect 172480 147568 172486 147580
rect 193950 147568 193956 147580
rect 194008 147568 194014 147620
rect 171502 147500 171508 147552
rect 171560 147540 171566 147552
rect 176102 147540 176108 147552
rect 171560 147512 176108 147540
rect 171560 147500 171566 147512
rect 176102 147500 176108 147512
rect 176160 147500 176166 147552
rect 371326 147228 371332 147280
rect 371384 147268 371390 147280
rect 375558 147268 375564 147280
rect 371384 147240 375564 147268
rect 371384 147228 371390 147240
rect 375558 147228 375564 147240
rect 375616 147228 375622 147280
rect 513374 147092 513380 147144
rect 513432 147132 513438 147144
rect 513558 147132 513564 147144
rect 513432 147104 513564 147132
rect 513432 147092 513438 147104
rect 513558 147092 513564 147104
rect 513616 147092 513622 147144
rect 513650 147024 513656 147076
rect 513708 147064 513714 147076
rect 514478 147064 514484 147076
rect 513708 147036 514484 147064
rect 513708 147024 513714 147036
rect 514478 147024 514484 147036
rect 514536 147024 514542 147076
rect 513558 146956 513564 147008
rect 513616 146996 513622 147008
rect 514386 146996 514392 147008
rect 513616 146968 514392 146996
rect 513616 146956 513622 146968
rect 514386 146956 514392 146968
rect 514444 146956 514450 147008
rect 513742 146888 513748 146940
rect 513800 146928 513806 146940
rect 514570 146928 514576 146940
rect 513800 146900 514576 146928
rect 513800 146888 513806 146900
rect 514570 146888 514576 146900
rect 514628 146888 514634 146940
rect 369210 146820 369216 146872
rect 369268 146860 369274 146872
rect 369762 146860 369768 146872
rect 369268 146832 369768 146860
rect 369268 146820 369274 146832
rect 369762 146820 369768 146832
rect 369820 146820 369826 146872
rect 371970 146820 371976 146872
rect 372028 146860 372034 146872
rect 375650 146860 375656 146872
rect 372028 146832 375656 146860
rect 372028 146820 372034 146832
rect 375650 146820 375656 146832
rect 375708 146820 375714 146872
rect 372614 146752 372620 146804
rect 372672 146792 372678 146804
rect 373718 146792 373724 146804
rect 372672 146764 373724 146792
rect 372672 146752 372678 146764
rect 373718 146752 373724 146764
rect 373776 146752 373782 146804
rect 182910 146276 182916 146328
rect 182968 146316 182974 146328
rect 197630 146316 197636 146328
rect 182968 146288 197636 146316
rect 182968 146276 182974 146288
rect 197630 146276 197636 146288
rect 197688 146276 197694 146328
rect 172422 146208 172428 146260
rect 172480 146248 172486 146260
rect 196802 146248 196808 146260
rect 172480 146220 196808 146248
rect 172480 146208 172486 146220
rect 196802 146208 196808 146220
rect 196860 146208 196866 146260
rect 371970 146208 371976 146260
rect 372028 146248 372034 146260
rect 393958 146248 393964 146260
rect 372028 146220 393964 146248
rect 372028 146208 372034 146220
rect 393958 146208 393964 146220
rect 394016 146208 394022 146260
rect 172330 146140 172336 146192
rect 172388 146180 172394 146192
rect 174722 146180 174728 146192
rect 172388 146152 174728 146180
rect 172388 146140 172394 146152
rect 174722 146140 174728 146152
rect 174780 146140 174786 146192
rect 171502 145800 171508 145852
rect 171560 145840 171566 145852
rect 178862 145840 178868 145852
rect 171560 145812 178868 145840
rect 171560 145800 171566 145812
rect 178862 145800 178868 145812
rect 178920 145800 178926 145852
rect 371326 145596 371332 145648
rect 371384 145636 371390 145648
rect 375926 145636 375932 145648
rect 371384 145608 375932 145636
rect 371384 145596 371390 145608
rect 375926 145596 375932 145608
rect 375984 145596 375990 145648
rect 371326 145460 371332 145512
rect 371384 145500 371390 145512
rect 375834 145500 375840 145512
rect 371384 145472 375840 145500
rect 371384 145460 371390 145472
rect 375834 145460 375840 145472
rect 375892 145460 375898 145512
rect 181530 144916 181536 144968
rect 181588 144956 181594 144968
rect 197354 144956 197360 144968
rect 181588 144928 197360 144956
rect 181588 144916 181594 144928
rect 197354 144916 197360 144928
rect 197412 144916 197418 144968
rect 172422 144848 172428 144900
rect 172480 144888 172486 144900
rect 195422 144888 195428 144900
rect 172480 144860 195428 144888
rect 172480 144848 172486 144860
rect 195422 144848 195428 144860
rect 195480 144848 195486 144900
rect 302786 144848 302792 144900
rect 302844 144888 302850 144900
rect 359642 144888 359648 144900
rect 302844 144860 359648 144888
rect 302844 144848 302850 144860
rect 359642 144848 359648 144860
rect 359700 144848 359706 144900
rect 515398 144848 515404 144900
rect 515456 144888 515462 144900
rect 516134 144888 516140 144900
rect 515456 144860 516140 144888
rect 515456 144848 515462 144860
rect 516134 144848 516140 144860
rect 516192 144848 516198 144900
rect 371326 144508 371332 144560
rect 371384 144548 371390 144560
rect 375742 144548 375748 144560
rect 371384 144520 375748 144548
rect 371384 144508 371390 144520
rect 375742 144508 375748 144520
rect 375800 144508 375806 144560
rect 171594 144168 171600 144220
rect 171652 144208 171658 144220
rect 184198 144208 184204 144220
rect 171652 144180 184204 144208
rect 171652 144168 171658 144180
rect 184198 144168 184204 144180
rect 184256 144168 184262 144220
rect 371326 144100 371332 144152
rect 371384 144140 371390 144152
rect 374454 144140 374460 144152
rect 371384 144112 374460 144140
rect 371384 144100 371390 144112
rect 374454 144100 374460 144112
rect 374512 144100 374518 144152
rect 172238 143488 172244 143540
rect 172296 143528 172302 143540
rect 186958 143528 186964 143540
rect 172296 143500 186964 143528
rect 172296 143488 172302 143500
rect 186958 143488 186964 143500
rect 187016 143488 187022 143540
rect 406378 143528 406384 143540
rect 393286 143500 406384 143528
rect 371326 143420 371332 143472
rect 371384 143460 371390 143472
rect 393286 143460 393314 143500
rect 406378 143488 406384 143500
rect 406436 143528 406442 143540
rect 431402 143528 431408 143540
rect 406436 143500 431408 143528
rect 406436 143488 406442 143500
rect 431402 143488 431408 143500
rect 431460 143488 431466 143540
rect 371384 143432 393314 143460
rect 371384 143420 371390 143432
rect 371970 143012 371976 143064
rect 372028 143052 372034 143064
rect 372982 143052 372988 143064
rect 372028 143024 372988 143052
rect 372028 143012 372034 143024
rect 372982 143012 372988 143024
rect 373040 143012 373046 143064
rect 171502 142808 171508 142860
rect 171560 142848 171566 142860
rect 182818 142848 182824 142860
rect 171560 142820 182824 142848
rect 171560 142808 171566 142820
rect 182818 142808 182824 142820
rect 182876 142808 182882 142860
rect 179414 142128 179420 142180
rect 179472 142168 179478 142180
rect 197354 142168 197360 142180
rect 179472 142140 197360 142168
rect 179472 142128 179478 142140
rect 197354 142128 197360 142140
rect 197412 142128 197418 142180
rect 172422 142060 172428 142112
rect 172480 142100 172486 142112
rect 181438 142100 181444 142112
rect 172480 142072 181444 142100
rect 172480 142060 172486 142072
rect 181438 142060 181444 142072
rect 181496 142060 181502 142112
rect 302326 142060 302332 142112
rect 302384 142100 302390 142112
rect 359550 142100 359556 142112
rect 302384 142072 359556 142100
rect 302384 142060 302390 142072
rect 359550 142060 359556 142072
rect 359608 142060 359614 142112
rect 371970 142060 371976 142112
rect 372028 142100 372034 142112
rect 381538 142100 381544 142112
rect 372028 142072 381544 142100
rect 372028 142060 372034 142072
rect 381538 142060 381544 142072
rect 381596 142100 381602 142112
rect 431310 142100 431316 142112
rect 381596 142072 431316 142100
rect 381596 142060 381602 142072
rect 431310 142060 431316 142072
rect 431368 142060 431374 142112
rect 171410 141924 171416 141976
rect 171468 141964 171474 141976
rect 178770 141964 178776 141976
rect 171468 141936 178776 141964
rect 171468 141924 171474 141936
rect 178770 141924 178776 141936
rect 178828 141924 178834 141976
rect 171502 141244 171508 141296
rect 171560 141284 171566 141296
rect 180058 141284 180064 141296
rect 171560 141256 180064 141284
rect 171560 141244 171566 141256
rect 180058 141244 180064 141256
rect 180116 141244 180122 141296
rect 178034 140768 178040 140820
rect 178092 140808 178098 140820
rect 197354 140808 197360 140820
rect 178092 140780 197360 140808
rect 178092 140768 178098 140780
rect 197354 140768 197360 140780
rect 197412 140768 197418 140820
rect 372614 140360 372620 140412
rect 372672 140400 372678 140412
rect 372982 140400 372988 140412
rect 372672 140372 372988 140400
rect 372672 140360 372678 140372
rect 372982 140360 372988 140372
rect 373040 140360 373046 140412
rect 172238 140020 172244 140072
rect 172296 140060 172302 140072
rect 187050 140060 187056 140072
rect 172296 140032 187056 140060
rect 172296 140020 172302 140032
rect 187050 140020 187056 140032
rect 187108 140020 187114 140072
rect 171686 139748 171692 139800
rect 171744 139788 171750 139800
rect 173158 139788 173164 139800
rect 171744 139760 173164 139788
rect 171744 139748 171750 139760
rect 173158 139748 173164 139760
rect 173216 139748 173222 139800
rect 371694 139340 371700 139392
rect 371752 139380 371758 139392
rect 371970 139380 371976 139392
rect 371752 139352 371976 139380
rect 371752 139340 371758 139352
rect 371970 139340 371976 139352
rect 372028 139340 372034 139392
rect 372154 139340 372160 139392
rect 372212 139380 372218 139392
rect 372890 139380 372896 139392
rect 372212 139352 372896 139380
rect 372212 139340 372218 139352
rect 372890 139340 372896 139352
rect 372948 139340 372954 139392
rect 518158 139340 518164 139392
rect 518216 139380 518222 139392
rect 580166 139380 580172 139392
rect 518216 139352 580172 139380
rect 518216 139340 518222 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 172422 139272 172428 139324
rect 172480 139312 172486 139324
rect 177390 139312 177396 139324
rect 172480 139284 177396 139312
rect 172480 139272 172486 139284
rect 177390 139272 177396 139284
rect 177448 139272 177454 139324
rect 371326 139272 371332 139324
rect 371384 139312 371390 139324
rect 395338 139312 395344 139324
rect 371384 139284 395344 139312
rect 371384 139272 371390 139284
rect 395338 139272 395344 139284
rect 395396 139312 395402 139324
rect 395982 139312 395988 139324
rect 395396 139284 395988 139312
rect 395396 139272 395402 139284
rect 395982 139272 395988 139284
rect 396040 139272 396046 139324
rect 371694 139204 371700 139256
rect 371752 139244 371758 139256
rect 399478 139244 399484 139256
rect 371752 139216 399484 139244
rect 371752 139204 371758 139216
rect 399478 139204 399484 139216
rect 399536 139204 399542 139256
rect 171870 138864 171876 138916
rect 171928 138904 171934 138916
rect 175918 138904 175924 138916
rect 171928 138876 175924 138904
rect 171928 138864 171934 138876
rect 175918 138864 175924 138876
rect 175976 138864 175982 138916
rect 171686 138728 171692 138780
rect 171744 138768 171750 138780
rect 174538 138768 174544 138780
rect 171744 138740 174544 138768
rect 171744 138728 171750 138740
rect 174538 138728 174544 138740
rect 174596 138728 174602 138780
rect 399478 138728 399484 138780
rect 399536 138768 399542 138780
rect 431310 138768 431316 138780
rect 399536 138740 431316 138768
rect 399536 138728 399542 138740
rect 431310 138728 431316 138740
rect 431368 138728 431374 138780
rect 395982 138660 395988 138712
rect 396040 138700 396046 138712
rect 429838 138700 429844 138712
rect 396040 138672 429844 138700
rect 396040 138660 396046 138672
rect 429838 138660 429844 138672
rect 429896 138660 429902 138712
rect 175918 137980 175924 138032
rect 175976 138020 175982 138032
rect 197354 138020 197360 138032
rect 175976 137992 197360 138020
rect 175976 137980 175982 137992
rect 197354 137980 197360 137992
rect 197412 137980 197418 138032
rect 445846 137980 445852 138032
rect 445904 138020 445910 138032
rect 446398 138020 446404 138032
rect 445904 137992 446404 138020
rect 445904 137980 445910 137992
rect 446398 137980 446404 137992
rect 446456 137980 446462 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 152458 137952 152464 137964
rect 3292 137924 152464 137952
rect 3292 137912 3298 137924
rect 152458 137912 152464 137924
rect 152516 137912 152522 137964
rect 172422 137912 172428 137964
rect 172480 137952 172486 137964
rect 188338 137952 188344 137964
rect 172480 137924 188344 137952
rect 172480 137912 172486 137924
rect 188338 137912 188344 137924
rect 188396 137912 188402 137964
rect 371326 137572 371332 137624
rect 371384 137612 371390 137624
rect 373626 137612 373632 137624
rect 371384 137584 373632 137612
rect 371384 137572 371390 137584
rect 373626 137572 373632 137584
rect 373684 137572 373690 137624
rect 371326 137300 371332 137352
rect 371384 137340 371390 137352
rect 371510 137340 371516 137352
rect 371384 137312 371516 137340
rect 371384 137300 371390 137312
rect 371510 137300 371516 137312
rect 371568 137300 371574 137352
rect 172330 137232 172336 137284
rect 172388 137272 172394 137284
rect 184290 137272 184296 137284
rect 172388 137244 184296 137272
rect 172388 137232 172394 137244
rect 184290 137232 184296 137244
rect 184348 137232 184354 137284
rect 172514 136620 172520 136672
rect 172572 136660 172578 136672
rect 197354 136660 197360 136672
rect 172572 136632 197360 136660
rect 172572 136620 172578 136632
rect 197354 136620 197360 136632
rect 197412 136620 197418 136672
rect 445294 136620 445300 136672
rect 445352 136660 445358 136672
rect 497458 136660 497464 136672
rect 445352 136632 497464 136660
rect 445352 136620 445358 136632
rect 497458 136620 497464 136632
rect 497516 136620 497522 136672
rect 172422 136552 172428 136604
rect 172480 136592 172486 136604
rect 182910 136592 182916 136604
rect 172480 136564 182916 136592
rect 172480 136552 172486 136564
rect 182910 136552 182916 136564
rect 182968 136552 182974 136604
rect 172238 136484 172244 136536
rect 172296 136524 172302 136536
rect 181530 136524 181536 136536
rect 172296 136496 181536 136524
rect 172296 136484 172302 136496
rect 181530 136484 181536 136496
rect 181588 136484 181594 136536
rect 170398 135872 170404 135924
rect 170456 135912 170462 135924
rect 197998 135912 198004 135924
rect 170456 135884 198004 135912
rect 170456 135872 170462 135884
rect 197998 135872 198004 135884
rect 198056 135872 198062 135924
rect 441614 135872 441620 135924
rect 441672 135912 441678 135924
rect 447226 135912 447232 135924
rect 441672 135884 447232 135912
rect 441672 135872 441678 135884
rect 447226 135872 447232 135884
rect 447284 135912 447290 135924
rect 500218 135912 500224 135924
rect 447284 135884 500224 135912
rect 447284 135872 447290 135884
rect 500218 135872 500224 135884
rect 500276 135872 500282 135924
rect 172238 135260 172244 135312
rect 172296 135300 172302 135312
rect 179414 135300 179420 135312
rect 172296 135272 179420 135300
rect 172296 135260 172302 135272
rect 179414 135260 179420 135272
rect 179472 135260 179478 135312
rect 445018 135260 445024 135312
rect 445076 135300 445082 135312
rect 445662 135300 445668 135312
rect 445076 135272 445668 135300
rect 445076 135260 445082 135272
rect 445662 135260 445668 135272
rect 445720 135300 445726 135312
rect 503070 135300 503076 135312
rect 445720 135272 503076 135300
rect 445720 135260 445726 135272
rect 503070 135260 503076 135272
rect 503128 135260 503134 135312
rect 171686 135192 171692 135244
rect 171744 135232 171750 135244
rect 175918 135232 175924 135244
rect 171744 135204 175924 135232
rect 171744 135192 171750 135204
rect 175918 135192 175924 135204
rect 175976 135192 175982 135244
rect 369118 135192 369124 135244
rect 369176 135192 369182 135244
rect 171870 135124 171876 135176
rect 171928 135164 171934 135176
rect 178034 135164 178040 135176
rect 171928 135136 178040 135164
rect 171928 135124 171934 135136
rect 178034 135124 178040 135136
rect 178092 135124 178098 135176
rect 369136 134904 369164 135192
rect 369118 134852 369124 134904
rect 369176 134852 369182 134904
rect 371694 134308 371700 134360
rect 371752 134348 371758 134360
rect 374178 134348 374184 134360
rect 371752 134320 374184 134348
rect 371752 134308 371758 134320
rect 374178 134308 374184 134320
rect 374236 134308 374242 134360
rect 443086 133968 443092 134020
rect 443144 134008 443150 134020
rect 490558 134008 490564 134020
rect 443144 133980 490564 134008
rect 443144 133968 443150 133980
rect 490558 133968 490564 133980
rect 490616 133968 490622 134020
rect 172422 133900 172428 133952
rect 172480 133940 172486 133952
rect 197722 133940 197728 133952
rect 172480 133912 197728 133940
rect 172480 133900 172486 133912
rect 197722 133900 197728 133912
rect 197780 133900 197786 133952
rect 442902 133900 442908 133952
rect 442960 133940 442966 133952
rect 445110 133940 445116 133952
rect 442960 133912 445116 133940
rect 442960 133900 442966 133912
rect 445110 133900 445116 133912
rect 445168 133940 445174 133952
rect 503162 133940 503168 133952
rect 445168 133912 503168 133940
rect 445168 133900 445174 133912
rect 503162 133900 503168 133912
rect 503220 133900 503226 133952
rect 371510 132948 371516 133000
rect 371568 132988 371574 133000
rect 372982 132988 372988 133000
rect 371568 132960 372988 132988
rect 371568 132948 371574 132960
rect 372982 132948 372988 132960
rect 373040 132948 373046 133000
rect 171134 132472 171140 132524
rect 171192 132512 171198 132524
rect 197354 132512 197360 132524
rect 171192 132484 197360 132512
rect 171192 132472 171198 132484
rect 197354 132472 197360 132484
rect 197412 132472 197418 132524
rect 442810 132472 442816 132524
rect 442868 132512 442874 132524
rect 444190 132512 444196 132524
rect 442868 132484 444196 132512
rect 442868 132472 442874 132484
rect 444190 132472 444196 132484
rect 444248 132472 444254 132524
rect 445110 132472 445116 132524
rect 445168 132512 445174 132524
rect 503254 132512 503260 132524
rect 445168 132484 503260 132512
rect 445168 132472 445174 132484
rect 503254 132472 503260 132484
rect 503312 132472 503318 132524
rect 172422 131044 172428 131096
rect 172480 131084 172486 131096
rect 197354 131084 197360 131096
rect 172480 131056 197360 131084
rect 172480 131044 172486 131056
rect 197354 131044 197360 131056
rect 197412 131044 197418 131096
rect 370038 130432 370044 130484
rect 370096 130472 370102 130484
rect 373258 130472 373264 130484
rect 370096 130444 373264 130472
rect 370096 130432 370102 130444
rect 373258 130432 373264 130444
rect 373316 130432 373322 130484
rect 370314 130364 370320 130416
rect 370372 130404 370378 130416
rect 373350 130404 373356 130416
rect 370372 130376 373356 130404
rect 370372 130364 370378 130376
rect 373350 130364 373356 130376
rect 373408 130364 373414 130416
rect 172238 129956 172244 130008
rect 172296 129996 172302 130008
rect 178034 129996 178040 130008
rect 172296 129968 178040 129996
rect 172296 129956 172302 129968
rect 178034 129956 178040 129968
rect 178092 129956 178098 130008
rect 444834 129004 444840 129056
rect 444892 129044 444898 129056
rect 476758 129044 476764 129056
rect 444892 129016 476764 129044
rect 444892 129004 444898 129016
rect 476758 129004 476764 129016
rect 476816 129044 476822 129056
rect 503622 129044 503628 129056
rect 476816 129016 503628 129044
rect 476816 129004 476822 129016
rect 503622 129004 503628 129016
rect 503680 129004 503686 129056
rect 172330 128256 172336 128308
rect 172388 128296 172394 128308
rect 197354 128296 197360 128308
rect 172388 128268 197360 128296
rect 172388 128256 172394 128268
rect 197354 128256 197360 128268
rect 197412 128256 197418 128308
rect 442902 127644 442908 127696
rect 442960 127684 442966 127696
rect 504266 127684 504272 127696
rect 442960 127656 504272 127684
rect 442960 127644 442966 127656
rect 504266 127644 504272 127656
rect 504324 127644 504330 127696
rect 443362 127576 443368 127628
rect 443420 127616 443426 127628
rect 444926 127616 444932 127628
rect 443420 127588 444932 127616
rect 443420 127576 443426 127588
rect 444926 127576 444932 127588
rect 444984 127616 444990 127628
rect 504358 127616 504364 127628
rect 444984 127588 504364 127616
rect 444984 127576 444990 127588
rect 504358 127576 504364 127588
rect 504416 127576 504422 127628
rect 171318 126896 171324 126948
rect 171376 126936 171382 126948
rect 197630 126936 197636 126948
rect 171376 126908 197636 126936
rect 171376 126896 171382 126908
rect 197630 126896 197636 126908
rect 197688 126896 197694 126948
rect 526438 126896 526444 126948
rect 526496 126936 526502 126948
rect 580166 126936 580172 126948
rect 526496 126908 580172 126936
rect 526496 126896 526502 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 444926 126284 444932 126336
rect 444984 126324 444990 126336
rect 467098 126324 467104 126336
rect 444984 126296 467104 126324
rect 444984 126284 444990 126296
rect 467098 126284 467104 126296
rect 467156 126324 467162 126336
rect 493962 126324 493968 126336
rect 467156 126296 493968 126324
rect 467156 126284 467162 126296
rect 493962 126284 493968 126296
rect 494020 126284 494026 126336
rect 444834 126216 444840 126268
rect 444892 126256 444898 126268
rect 457438 126256 457444 126268
rect 444892 126228 457444 126256
rect 444892 126216 444898 126228
rect 457438 126216 457444 126228
rect 457496 126256 457502 126268
rect 494698 126256 494704 126268
rect 457496 126228 494704 126256
rect 457496 126216 457502 126228
rect 494698 126216 494704 126228
rect 494756 126216 494762 126268
rect 371602 126012 371608 126064
rect 371660 126052 371666 126064
rect 441890 126052 441896 126064
rect 371660 126024 441896 126052
rect 371660 126012 371666 126024
rect 441890 126012 441896 126024
rect 441948 126012 441954 126064
rect 371694 125944 371700 125996
rect 371752 125984 371758 125996
rect 442902 125984 442908 125996
rect 371752 125956 442908 125984
rect 371752 125944 371758 125956
rect 442902 125944 442908 125956
rect 442960 125944 442966 125996
rect 370406 125876 370412 125928
rect 370464 125916 370470 125928
rect 371326 125916 371332 125928
rect 370464 125888 371332 125916
rect 370464 125876 370470 125888
rect 371326 125876 371332 125888
rect 371384 125916 371390 125928
rect 443362 125916 443368 125928
rect 371384 125888 443368 125916
rect 371384 125876 371390 125888
rect 443362 125876 443368 125888
rect 443420 125876 443426 125928
rect 172238 125740 172244 125792
rect 172296 125780 172302 125792
rect 180058 125780 180064 125792
rect 172296 125752 180064 125780
rect 172296 125740 172302 125752
rect 180058 125740 180064 125752
rect 180116 125740 180122 125792
rect 172422 125672 172428 125724
rect 172480 125712 172486 125724
rect 181438 125712 181444 125724
rect 172480 125684 181444 125712
rect 172480 125672 172486 125684
rect 181438 125672 181444 125684
rect 181496 125672 181502 125724
rect 172330 125604 172336 125656
rect 172388 125644 172394 125656
rect 182818 125644 182824 125656
rect 172388 125616 182824 125644
rect 172388 125604 172394 125616
rect 182818 125604 182824 125616
rect 182876 125604 182882 125656
rect 371418 125468 371424 125520
rect 371476 125508 371482 125520
rect 441798 125508 441804 125520
rect 371476 125480 441804 125508
rect 371476 125468 371482 125480
rect 441798 125468 441804 125480
rect 441856 125508 441862 125520
rect 444926 125508 444932 125520
rect 441856 125480 444932 125508
rect 441856 125468 441862 125480
rect 444926 125468 444932 125480
rect 444984 125468 444990 125520
rect 369302 125400 369308 125452
rect 369360 125440 369366 125452
rect 443086 125440 443092 125452
rect 369360 125412 443092 125440
rect 369360 125400 369366 125412
rect 443086 125400 443092 125412
rect 443144 125400 443150 125452
rect 374822 125332 374828 125384
rect 374880 125372 374886 125384
rect 442074 125372 442080 125384
rect 374880 125344 442080 125372
rect 374880 125332 374886 125344
rect 442074 125332 442080 125344
rect 442132 125372 442138 125384
rect 444834 125372 444840 125384
rect 442132 125344 444840 125372
rect 442132 125332 442138 125344
rect 444834 125332 444840 125344
rect 444892 125332 444898 125384
rect 441614 125304 441620 125316
rect 373966 125276 441620 125304
rect 302418 125196 302424 125248
rect 302476 125236 302482 125248
rect 369946 125236 369952 125248
rect 302476 125208 369952 125236
rect 302476 125196 302482 125208
rect 369946 125196 369952 125208
rect 370004 125196 370010 125248
rect 302510 125128 302516 125180
rect 302568 125168 302574 125180
rect 369854 125168 369860 125180
rect 302568 125140 369860 125168
rect 302568 125128 302574 125140
rect 369854 125128 369860 125140
rect 369912 125168 369918 125180
rect 373966 125168 373994 125276
rect 441614 125264 441620 125276
rect 441672 125264 441678 125316
rect 445754 125236 445760 125248
rect 369912 125140 373994 125168
rect 441586 125208 445760 125236
rect 369912 125128 369918 125140
rect 302878 125060 302884 125112
rect 302936 125100 302942 125112
rect 370038 125100 370044 125112
rect 302936 125072 370044 125100
rect 302936 125060 302942 125072
rect 370038 125060 370044 125072
rect 370096 125060 370102 125112
rect 302694 124992 302700 125044
rect 302752 125032 302758 125044
rect 369302 125032 369308 125044
rect 302752 125004 369308 125032
rect 302752 124992 302758 125004
rect 369302 124992 369308 125004
rect 369360 124992 369366 125044
rect 302970 124924 302976 124976
rect 303028 124964 303034 124976
rect 370314 124964 370320 124976
rect 303028 124936 370320 124964
rect 303028 124924 303034 124936
rect 370314 124924 370320 124936
rect 370372 124924 370378 124976
rect 441586 124908 441614 125208
rect 445754 125196 445760 125208
rect 445812 125236 445818 125248
rect 513190 125236 513196 125248
rect 445812 125208 513196 125236
rect 445812 125196 445818 125208
rect 513190 125196 513196 125208
rect 513248 125196 513254 125248
rect 493962 125128 493968 125180
rect 494020 125168 494026 125180
rect 513374 125168 513380 125180
rect 494020 125140 513380 125168
rect 494020 125128 494026 125140
rect 513374 125128 513380 125140
rect 513432 125128 513438 125180
rect 494698 125060 494704 125112
rect 494756 125100 494762 125112
rect 494756 125072 513420 125100
rect 494756 125060 494762 125072
rect 513392 125044 513420 125072
rect 500218 124992 500224 125044
rect 500276 125032 500282 125044
rect 513282 125032 513288 125044
rect 500276 125004 513288 125032
rect 500276 124992 500282 125004
rect 513282 124992 513288 125004
rect 513340 124992 513346 125044
rect 513374 124992 513380 125044
rect 513432 124992 513438 125044
rect 446398 124924 446404 124976
rect 446456 124964 446462 124976
rect 516134 124964 516140 124976
rect 446456 124936 516140 124964
rect 446456 124924 446462 124936
rect 516134 124924 516140 124936
rect 516192 124924 516198 124976
rect 172514 124856 172520 124908
rect 172572 124896 172578 124908
rect 197446 124896 197452 124908
rect 172572 124868 197452 124896
rect 172572 124856 172578 124868
rect 197446 124856 197452 124868
rect 197504 124856 197510 124908
rect 302234 124856 302240 124908
rect 302292 124896 302298 124908
rect 370222 124896 370228 124908
rect 302292 124868 370228 124896
rect 302292 124856 302298 124868
rect 370222 124856 370228 124868
rect 370280 124856 370286 124908
rect 370866 124856 370872 124908
rect 370924 124896 370930 124908
rect 441586 124896 441620 124908
rect 370924 124868 441620 124896
rect 370924 124856 370930 124868
rect 441614 124856 441620 124868
rect 441672 124856 441678 124908
rect 490558 124856 490564 124908
rect 490616 124896 490622 124908
rect 513466 124896 513472 124908
rect 490616 124868 513472 124896
rect 490616 124856 490622 124868
rect 513466 124856 513472 124868
rect 513524 124856 513530 124908
rect 497458 124788 497464 124840
rect 497516 124828 497522 124840
rect 516226 124828 516232 124840
rect 497516 124800 516232 124828
rect 497516 124788 497522 124800
rect 516226 124788 516232 124800
rect 516284 124788 516290 124840
rect 369854 124720 369860 124772
rect 369912 124760 369918 124772
rect 374086 124760 374092 124772
rect 369912 124732 374092 124760
rect 369912 124720 369918 124732
rect 374086 124720 374092 124732
rect 374144 124760 374150 124772
rect 374822 124760 374828 124772
rect 374144 124732 374828 124760
rect 374144 124720 374150 124732
rect 374822 124720 374828 124732
rect 374880 124720 374886 124772
rect 429838 124720 429844 124772
rect 429896 124760 429902 124772
rect 516318 124760 516324 124772
rect 429896 124732 516324 124760
rect 429896 124720 429902 124732
rect 516318 124720 516324 124732
rect 516376 124720 516382 124772
rect 171502 124312 171508 124364
rect 171560 124352 171566 124364
rect 175918 124352 175924 124364
rect 171560 124324 175924 124352
rect 171560 124312 171566 124324
rect 175918 124312 175924 124324
rect 175976 124312 175982 124364
rect 171870 124244 171876 124296
rect 171928 124284 171934 124296
rect 174538 124284 174544 124296
rect 171928 124256 174544 124284
rect 171928 124244 171934 124256
rect 174538 124244 174544 124256
rect 174596 124244 174602 124296
rect 172146 124176 172152 124228
rect 172204 124216 172210 124228
rect 173158 124216 173164 124228
rect 172204 124188 173164 124216
rect 172204 124176 172210 124188
rect 173158 124176 173164 124188
rect 173216 124176 173222 124228
rect 178034 124108 178040 124160
rect 178092 124148 178098 124160
rect 197354 124148 197360 124160
rect 178092 124120 197360 124148
rect 178092 124108 178098 124120
rect 197354 124108 197360 124120
rect 197412 124108 197418 124160
rect 431310 124108 431316 124160
rect 431368 124148 431374 124160
rect 516502 124148 516508 124160
rect 431368 124120 516508 124148
rect 431368 124108 431374 124120
rect 516502 124108 516508 124120
rect 516560 124108 516566 124160
rect 368198 124040 368204 124092
rect 368256 124080 368262 124092
rect 369394 124080 369400 124092
rect 368256 124052 369400 124080
rect 368256 124040 368262 124052
rect 369394 124040 369400 124052
rect 369452 124040 369458 124092
rect 503070 124040 503076 124092
rect 503128 124080 503134 124092
rect 513834 124080 513840 124092
rect 503128 124052 513840 124080
rect 503128 124040 503134 124052
rect 513834 124040 513840 124052
rect 513892 124040 513898 124092
rect 503162 123972 503168 124024
rect 503220 124012 503226 124024
rect 513742 124012 513748 124024
rect 503220 123984 513748 124012
rect 503220 123972 503226 123984
rect 513742 123972 513748 123984
rect 513800 123972 513806 124024
rect 503622 123904 503628 123956
rect 503680 123944 503686 123956
rect 513558 123944 513564 123956
rect 503680 123916 513564 123944
rect 503680 123904 503686 123916
rect 513558 123904 513564 123916
rect 513616 123904 513622 123956
rect 503254 123836 503260 123888
rect 503312 123876 503318 123888
rect 513926 123876 513932 123888
rect 503312 123848 513932 123876
rect 503312 123836 503318 123848
rect 513926 123836 513932 123848
rect 513984 123836 513990 123888
rect 504358 123768 504364 123820
rect 504416 123808 504422 123820
rect 513650 123808 513656 123820
rect 504416 123780 513656 123808
rect 504416 123768 504422 123780
rect 513650 123768 513656 123780
rect 513708 123768 513714 123820
rect 504266 123700 504272 123752
rect 504324 123740 504330 123752
rect 514110 123740 514116 123752
rect 504324 123712 514116 123740
rect 504324 123700 504330 123712
rect 514110 123700 514116 123712
rect 514168 123700 514174 123752
rect 302970 123496 302976 123548
rect 303028 123536 303034 123548
rect 370406 123536 370412 123548
rect 303028 123508 370412 123536
rect 303028 123496 303034 123508
rect 370406 123496 370412 123508
rect 370464 123496 370470 123548
rect 302878 123428 302884 123480
rect 302936 123468 302942 123480
rect 369854 123468 369860 123480
rect 302936 123440 369860 123468
rect 302936 123428 302942 123440
rect 369854 123428 369860 123440
rect 369912 123428 369918 123480
rect 168926 122884 168932 122936
rect 168984 122924 168990 122936
rect 177298 122924 177304 122936
rect 168984 122896 177304 122924
rect 168984 122884 168990 122896
rect 177298 122884 177304 122896
rect 177356 122884 177362 122936
rect 160922 122816 160928 122868
rect 160980 122856 160986 122868
rect 192478 122856 192484 122868
rect 160980 122828 192484 122856
rect 160980 122816 160986 122828
rect 192478 122816 192484 122828
rect 192536 122816 192542 122868
rect 320818 122816 320824 122868
rect 320876 122856 320882 122868
rect 510890 122856 510896 122868
rect 320876 122828 510896 122856
rect 320876 122816 320882 122828
rect 510890 122816 510896 122828
rect 510948 122816 510954 122868
rect 164878 122748 164884 122800
rect 164936 122788 164942 122800
rect 170398 122788 170404 122800
rect 164936 122760 170404 122788
rect 164936 122748 164942 122760
rect 170398 122748 170404 122760
rect 170456 122748 170462 122800
rect 191098 122788 191104 122800
rect 171106 122760 191104 122788
rect 162854 122680 162860 122732
rect 162912 122720 162918 122732
rect 171106 122720 171134 122760
rect 191098 122748 191104 122760
rect 191156 122748 191162 122800
rect 431862 122748 431868 122800
rect 431920 122788 431926 122800
rect 434714 122788 434720 122800
rect 431920 122760 434720 122788
rect 431920 122748 431926 122760
rect 434714 122748 434720 122760
rect 434772 122748 434778 122800
rect 441246 122748 441252 122800
rect 441304 122788 441310 122800
rect 512914 122788 512920 122800
rect 441304 122760 512920 122788
rect 441304 122748 441310 122760
rect 512914 122748 512920 122760
rect 512972 122748 512978 122800
rect 162912 122692 171134 122720
rect 162912 122680 162918 122692
rect 433150 122680 433156 122732
rect 433208 122720 433214 122732
rect 504910 122720 504916 122732
rect 433208 122692 504916 122720
rect 433208 122680 433214 122692
rect 504910 122680 504916 122692
rect 504968 122680 504974 122732
rect 506842 122680 506848 122732
rect 506900 122720 506906 122732
rect 514018 122720 514024 122732
rect 506900 122692 514024 122720
rect 506900 122680 506906 122692
rect 514018 122680 514024 122692
rect 514076 122680 514082 122732
rect 437198 122612 437204 122664
rect 437256 122652 437262 122664
rect 441706 122652 441712 122664
rect 437256 122624 441712 122652
rect 437256 122612 437262 122624
rect 441706 122612 441712 122624
rect 441764 122652 441770 122664
rect 508866 122652 508872 122664
rect 441764 122624 508872 122652
rect 441764 122612 441770 122624
rect 508866 122612 508872 122624
rect 508924 122612 508930 122664
rect 309778 122544 309784 122596
rect 309836 122584 309842 122596
rect 438854 122584 438860 122596
rect 309836 122556 438860 122584
rect 309836 122544 309842 122556
rect 438854 122544 438860 122556
rect 438912 122544 438918 122596
rect 301498 122068 301504 122120
rect 301556 122108 301562 122120
rect 366910 122108 366916 122120
rect 301556 122080 366916 122108
rect 301556 122068 301562 122080
rect 366910 122068 366916 122080
rect 366968 122068 366974 122120
rect 172054 120028 172060 120080
rect 172112 120068 172118 120080
rect 197354 120068 197360 120080
rect 172112 120040 197360 120068
rect 172112 120028 172118 120040
rect 197354 120028 197360 120040
rect 197412 120028 197418 120080
rect 302510 120028 302516 120080
rect 302568 120068 302574 120080
rect 370130 120068 370136 120080
rect 302568 120040 370136 120068
rect 302568 120028 302574 120040
rect 370130 120028 370136 120040
rect 370188 120028 370194 120080
rect 171870 118600 171876 118652
rect 171928 118640 171934 118652
rect 197630 118640 197636 118652
rect 171928 118612 197636 118640
rect 171928 118600 171934 118612
rect 197630 118600 197636 118612
rect 197688 118600 197694 118652
rect 302602 117240 302608 117292
rect 302660 117280 302666 117292
rect 368198 117280 368204 117292
rect 302660 117252 368204 117280
rect 302660 117240 302666 117252
rect 368198 117240 368204 117252
rect 368256 117240 368262 117292
rect 171962 115880 171968 115932
rect 172020 115920 172026 115932
rect 198550 115920 198556 115932
rect 172020 115892 198556 115920
rect 172020 115880 172026 115892
rect 198550 115880 198556 115892
rect 198608 115880 198614 115932
rect 171778 114452 171784 114504
rect 171836 114492 171842 114504
rect 197538 114492 197544 114504
rect 171836 114464 197544 114492
rect 171836 114452 171842 114464
rect 197538 114452 197544 114464
rect 197596 114452 197602 114504
rect 318058 113092 318064 113144
rect 318116 113132 318122 113144
rect 579798 113132 579804 113144
rect 318116 113104 579804 113132
rect 318116 113092 318122 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 175918 112412 175924 112464
rect 175976 112452 175982 112464
rect 197446 112452 197452 112464
rect 175976 112424 197452 112452
rect 175976 112412 175982 112424
rect 197446 112412 197452 112424
rect 197504 112412 197510 112464
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 159358 111772 159364 111784
rect 3476 111744 159364 111772
rect 3476 111732 3482 111744
rect 159358 111732 159364 111744
rect 159416 111732 159422 111784
rect 182818 111732 182824 111784
rect 182876 111772 182882 111784
rect 197354 111772 197360 111784
rect 182876 111744 197360 111772
rect 182876 111732 182882 111744
rect 197354 111732 197360 111744
rect 197412 111732 197418 111784
rect 302510 111732 302516 111784
rect 302568 111772 302574 111784
rect 370498 111772 370504 111784
rect 302568 111744 370504 111772
rect 302568 111732 302574 111744
rect 370498 111732 370504 111744
rect 370556 111732 370562 111784
rect 181438 110372 181444 110424
rect 181496 110412 181502 110424
rect 197538 110412 197544 110424
rect 181496 110384 197544 110412
rect 181496 110372 181502 110384
rect 197538 110372 197544 110384
rect 197596 110372 197602 110424
rect 302786 108944 302792 108996
rect 302844 108984 302850 108996
rect 371418 108984 371424 108996
rect 302844 108956 371424 108984
rect 302844 108944 302850 108956
rect 371418 108944 371424 108956
rect 371476 108944 371482 108996
rect 180058 107584 180064 107636
rect 180116 107624 180122 107636
rect 197998 107624 198004 107636
rect 180116 107596 198004 107624
rect 180116 107584 180122 107596
rect 197998 107584 198004 107596
rect 198056 107584 198062 107636
rect 174538 103436 174544 103488
rect 174596 103476 174602 103488
rect 197998 103476 198004 103488
rect 174596 103448 198004 103476
rect 174596 103436 174602 103448
rect 197998 103436 198004 103448
rect 198056 103436 198062 103488
rect 173158 102076 173164 102128
rect 173216 102116 173222 102128
rect 197998 102116 198004 102128
rect 173216 102088 198004 102116
rect 173216 102076 173222 102088
rect 197998 102076 198004 102088
rect 198056 102076 198062 102128
rect 302786 102076 302792 102128
rect 302844 102116 302850 102128
rect 369854 102116 369860 102128
rect 302844 102088 369860 102116
rect 302844 102076 302850 102088
rect 369854 102076 369860 102088
rect 369912 102076 369918 102128
rect 533338 100648 533344 100700
rect 533396 100688 533402 100700
rect 580166 100688 580172 100700
rect 533396 100660 580172 100688
rect 533396 100648 533402 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 232038 99968 232044 100020
rect 232096 100008 232102 100020
rect 232096 99980 232360 100008
rect 232096 99968 232102 99980
rect 232332 99952 232360 99980
rect 232314 99900 232320 99952
rect 232372 99900 232378 99952
rect 298922 99696 298928 99748
rect 298980 99736 298986 99748
rect 322198 99736 322204 99748
rect 298980 99708 322204 99736
rect 298980 99696 298986 99708
rect 322198 99696 322204 99708
rect 322256 99696 322262 99748
rect 299106 99628 299112 99680
rect 299164 99668 299170 99680
rect 323578 99668 323584 99680
rect 299164 99640 323584 99668
rect 299164 99628 299170 99640
rect 323578 99628 323584 99640
rect 323636 99628 323642 99680
rect 298646 99560 298652 99612
rect 298704 99600 298710 99612
rect 359458 99600 359464 99612
rect 298704 99572 359464 99600
rect 298704 99560 298710 99572
rect 359458 99560 359464 99572
rect 359516 99560 359522 99612
rect 299474 99492 299480 99544
rect 299532 99532 299538 99544
rect 431218 99532 431224 99544
rect 299532 99504 431224 99532
rect 299532 99492 299538 99504
rect 431218 99492 431224 99504
rect 431276 99492 431282 99544
rect 211614 99424 211620 99476
rect 211672 99464 211678 99476
rect 211798 99464 211804 99476
rect 211672 99436 211804 99464
rect 211672 99424 211678 99436
rect 211798 99424 211804 99436
rect 211856 99424 211862 99476
rect 299842 99424 299848 99476
rect 299900 99464 299906 99476
rect 501598 99464 501604 99476
rect 299900 99436 501604 99464
rect 299900 99424 299906 99436
rect 501598 99424 501604 99436
rect 501656 99424 501662 99476
rect 166902 99356 166908 99408
rect 166960 99396 166966 99408
rect 298278 99396 298284 99408
rect 166960 99368 298284 99396
rect 166960 99356 166966 99368
rect 298278 99356 298284 99368
rect 298336 99356 298342 99408
rect 299658 99356 299664 99408
rect 299716 99396 299722 99408
rect 502978 99396 502984 99408
rect 299716 99368 502984 99396
rect 299716 99356 299722 99368
rect 502978 99356 502984 99368
rect 503036 99356 503042 99408
rect 298462 99288 298468 99340
rect 298520 99328 298526 99340
rect 301498 99328 301504 99340
rect 298520 99300 301504 99328
rect 298520 99288 298526 99300
rect 301498 99288 301504 99300
rect 301556 99288 301562 99340
rect 305730 99328 305736 99340
rect 302206 99300 305736 99328
rect 101398 99220 101404 99272
rect 101456 99260 101462 99272
rect 211982 99260 211988 99272
rect 101456 99232 211988 99260
rect 101456 99220 101462 99232
rect 211982 99220 211988 99232
rect 212040 99220 212046 99272
rect 299290 99220 299296 99272
rect 299348 99260 299354 99272
rect 302206 99260 302234 99300
rect 305730 99288 305736 99300
rect 305788 99288 305794 99340
rect 299348 99232 302234 99260
rect 299348 99220 299354 99232
rect 94498 99152 94504 99204
rect 94556 99192 94562 99204
rect 207842 99192 207848 99204
rect 94556 99164 207848 99192
rect 94556 99152 94562 99164
rect 207842 99152 207848 99164
rect 207900 99152 207906 99204
rect 271414 99152 271420 99204
rect 271472 99192 271478 99204
rect 423766 99192 423772 99204
rect 271472 99164 423772 99192
rect 271472 99152 271478 99164
rect 423766 99152 423772 99164
rect 423824 99152 423830 99204
rect 93118 99084 93124 99136
rect 93176 99124 93182 99136
rect 213822 99124 213828 99136
rect 93176 99096 213828 99124
rect 93176 99084 93182 99096
rect 213822 99084 213828 99096
rect 213880 99084 213886 99136
rect 273806 99084 273812 99136
rect 273864 99124 273870 99136
rect 435358 99124 435364 99136
rect 273864 99096 435364 99124
rect 273864 99084 273870 99096
rect 435358 99084 435364 99096
rect 435416 99084 435422 99136
rect 71038 99016 71044 99068
rect 71096 99056 71102 99068
rect 210234 99056 210240 99068
rect 71096 99028 210240 99056
rect 71096 99016 71102 99028
rect 210234 99016 210240 99028
rect 210292 99016 210298 99068
rect 275002 99016 275008 99068
rect 275060 99056 275066 99068
rect 440878 99056 440884 99068
rect 275060 99028 440884 99056
rect 275060 99016 275066 99028
rect 440878 99016 440884 99028
rect 440936 99016 440942 99068
rect 57238 98948 57244 99000
rect 57296 98988 57302 99000
rect 207658 98988 207664 99000
rect 57296 98960 207664 98988
rect 57296 98948 57302 98960
rect 207658 98948 207664 98960
rect 207716 98948 207722 99000
rect 290090 98948 290096 99000
rect 290148 98988 290154 99000
rect 457438 98988 457444 99000
rect 290148 98960 457444 98988
rect 290148 98948 290154 98960
rect 457438 98948 457444 98960
rect 457496 98948 457502 99000
rect 50338 98880 50344 98932
rect 50396 98920 50402 98932
rect 207014 98920 207020 98932
rect 50396 98892 207020 98920
rect 50396 98880 50402 98892
rect 207014 98880 207020 98892
rect 207072 98880 207078 98932
rect 277394 98880 277400 98932
rect 277452 98920 277458 98932
rect 458174 98920 458180 98932
rect 277452 98892 458180 98920
rect 277452 98880 277458 98892
rect 458174 98880 458180 98892
rect 458232 98880 458238 98932
rect 46198 98812 46204 98864
rect 46256 98852 46262 98864
rect 205818 98852 205824 98864
rect 46256 98824 205824 98852
rect 46256 98812 46262 98824
rect 205818 98812 205824 98824
rect 205876 98812 205882 98864
rect 279142 98812 279148 98864
rect 279200 98852 279206 98864
rect 467098 98852 467104 98864
rect 279200 98824 467104 98852
rect 279200 98812 279206 98824
rect 467098 98812 467104 98824
rect 467156 98812 467162 98864
rect 36538 98744 36544 98796
rect 36596 98784 36602 98796
rect 202230 98784 202236 98796
rect 36596 98756 202236 98784
rect 36596 98744 36602 98756
rect 202230 98744 202236 98756
rect 202288 98744 202294 98796
rect 282914 98744 282920 98796
rect 282972 98784 282978 98796
rect 490558 98784 490564 98796
rect 282972 98756 490564 98784
rect 282972 98744 282978 98756
rect 490558 98744 490564 98756
rect 490616 98744 490622 98796
rect 29638 98676 29644 98728
rect 29696 98716 29702 98728
rect 204622 98716 204628 98728
rect 29696 98688 204628 98716
rect 29696 98676 29702 98688
rect 204622 98676 204628 98688
rect 204680 98676 204686 98728
rect 292942 98676 292948 98728
rect 293000 98716 293006 98728
rect 550634 98716 550640 98728
rect 293000 98688 550640 98716
rect 293000 98676 293006 98688
rect 550634 98676 550640 98688
rect 550692 98676 550698 98728
rect 19242 98608 19248 98660
rect 19300 98648 19306 98660
rect 203058 98648 203064 98660
rect 19300 98620 203064 98648
rect 19300 98608 19306 98620
rect 203058 98608 203064 98620
rect 203116 98608 203122 98660
rect 293494 98608 293500 98660
rect 293552 98648 293558 98660
rect 554774 98648 554780 98660
rect 293552 98620 554780 98648
rect 293552 98608 293558 98620
rect 554774 98608 554780 98620
rect 554832 98608 554838 98660
rect 263042 98540 263048 98592
rect 263100 98580 263106 98592
rect 373994 98580 374000 98592
rect 263100 98552 374000 98580
rect 263100 98540 263106 98552
rect 373994 98540 374000 98552
rect 374052 98540 374058 98592
rect 258626 98472 258632 98524
rect 258684 98512 258690 98524
rect 345658 98512 345664 98524
rect 258684 98484 345664 98512
rect 258684 98472 258690 98484
rect 345658 98472 345664 98484
rect 345716 98472 345722 98524
rect 256878 98404 256884 98456
rect 256936 98444 256942 98456
rect 335998 98444 336004 98456
rect 256936 98416 336004 98444
rect 256936 98404 256942 98416
rect 335998 98404 336004 98416
rect 336056 98404 336062 98456
rect 218514 98336 218520 98388
rect 218572 98376 218578 98388
rect 218974 98376 218980 98388
rect 218572 98348 218980 98376
rect 218572 98336 218578 98348
rect 218974 98336 218980 98348
rect 219032 98336 219038 98388
rect 270770 98336 270776 98388
rect 270828 98376 270834 98388
rect 413278 98376 413284 98388
rect 270828 98348 413284 98376
rect 270828 98336 270834 98348
rect 413278 98336 413284 98348
rect 413336 98336 413342 98388
rect 201586 98268 201592 98320
rect 201644 98308 201650 98320
rect 201862 98308 201868 98320
rect 201644 98280 201868 98308
rect 201644 98268 201650 98280
rect 201862 98268 201868 98280
rect 201920 98268 201926 98320
rect 208486 98268 208492 98320
rect 208544 98308 208550 98320
rect 208854 98308 208860 98320
rect 208544 98280 208860 98308
rect 208544 98268 208550 98280
rect 208854 98268 208860 98280
rect 208912 98268 208918 98320
rect 270954 98268 270960 98320
rect 271012 98308 271018 98320
rect 414658 98308 414664 98320
rect 271012 98280 414664 98308
rect 271012 98268 271018 98280
rect 414658 98268 414664 98280
rect 414716 98268 414722 98320
rect 289354 98200 289360 98252
rect 289412 98240 289418 98252
rect 289630 98240 289636 98252
rect 289412 98212 289636 98240
rect 289412 98200 289418 98212
rect 289630 98200 289636 98212
rect 289688 98200 289694 98252
rect 150342 97928 150348 97980
rect 150400 97968 150406 97980
rect 225138 97968 225144 97980
rect 150400 97940 225144 97968
rect 150400 97928 150406 97940
rect 225138 97928 225144 97940
rect 225196 97928 225202 97980
rect 238110 97928 238116 97980
rect 238168 97968 238174 97980
rect 238754 97968 238760 97980
rect 238168 97940 238760 97968
rect 238168 97928 238174 97940
rect 238754 97928 238760 97940
rect 238812 97928 238818 97980
rect 322198 97968 322204 97980
rect 272536 97940 322204 97968
rect 134518 97860 134524 97912
rect 134576 97900 134582 97912
rect 214374 97900 214380 97912
rect 134576 97872 214380 97900
rect 134576 97860 134582 97872
rect 214374 97860 214380 97872
rect 214432 97860 214438 97912
rect 215294 97860 215300 97912
rect 215352 97900 215358 97912
rect 222378 97900 222384 97912
rect 215352 97872 222384 97900
rect 215352 97860 215358 97872
rect 222378 97860 222384 97872
rect 222436 97860 222442 97912
rect 238018 97860 238024 97912
rect 238076 97900 238082 97912
rect 239674 97900 239680 97912
rect 238076 97872 239680 97900
rect 238076 97860 238082 97872
rect 239674 97860 239680 97872
rect 239732 97860 239738 97912
rect 126882 97792 126888 97844
rect 126940 97832 126946 97844
rect 126940 97804 210648 97832
rect 126940 97792 126946 97804
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 124858 97724 124864 97776
rect 124916 97764 124922 97776
rect 210620 97764 210648 97804
rect 215110 97792 215116 97844
rect 215168 97832 215174 97844
rect 219802 97832 219808 97844
rect 215168 97804 219808 97832
rect 215168 97792 215174 97804
rect 219802 97792 219808 97804
rect 219860 97792 219866 97844
rect 234614 97792 234620 97844
rect 234672 97832 234678 97844
rect 239306 97832 239312 97844
rect 234672 97804 239312 97832
rect 234672 97792 234678 97804
rect 239306 97792 239312 97804
rect 239364 97792 239370 97844
rect 251634 97792 251640 97844
rect 251692 97832 251698 97844
rect 256694 97832 256700 97844
rect 251692 97804 256700 97832
rect 251692 97792 251698 97804
rect 256694 97792 256700 97804
rect 256752 97792 256758 97844
rect 264606 97792 264612 97844
rect 264664 97832 264670 97844
rect 272536 97832 272564 97940
rect 322198 97928 322204 97940
rect 322256 97928 322262 97980
rect 272702 97860 272708 97912
rect 272760 97900 272766 97912
rect 327718 97900 327724 97912
rect 272760 97872 327724 97900
rect 272760 97860 272766 97872
rect 327718 97860 327724 97872
rect 327776 97860 327782 97912
rect 276014 97832 276020 97844
rect 264664 97804 272564 97832
rect 275296 97804 276020 97832
rect 264664 97792 264670 97804
rect 124916 97736 209084 97764
rect 210620 97736 215294 97764
rect 124916 97724 124922 97736
rect 126238 97656 126244 97708
rect 126296 97696 126302 97708
rect 208946 97696 208952 97708
rect 126296 97668 208952 97696
rect 126296 97656 126302 97668
rect 208946 97656 208952 97668
rect 209004 97656 209010 97708
rect 209056 97696 209084 97736
rect 215266 97696 215294 97736
rect 216674 97724 216680 97776
rect 216732 97764 216738 97776
rect 226334 97764 226340 97776
rect 216732 97736 226340 97764
rect 216732 97724 216738 97736
rect 226334 97724 226340 97736
rect 226392 97724 226398 97776
rect 242066 97724 242072 97776
rect 242124 97764 242130 97776
rect 253290 97764 253296 97776
rect 242124 97736 253296 97764
rect 242124 97724 242130 97736
rect 253290 97724 253296 97736
rect 253348 97724 253354 97776
rect 259270 97724 259276 97776
rect 259328 97764 259334 97776
rect 267274 97764 267280 97776
rect 259328 97736 267280 97764
rect 259328 97724 259334 97736
rect 267274 97724 267280 97736
rect 267332 97724 267338 97776
rect 268194 97724 268200 97776
rect 268252 97764 268258 97776
rect 275296 97764 275324 97804
rect 276014 97792 276020 97804
rect 276072 97792 276078 97844
rect 278130 97792 278136 97844
rect 278188 97832 278194 97844
rect 352558 97832 352564 97844
rect 278188 97804 352564 97832
rect 278188 97792 278194 97804
rect 352558 97792 352564 97804
rect 352616 97792 352622 97844
rect 268252 97736 275324 97764
rect 268252 97724 268258 97736
rect 275370 97724 275376 97776
rect 275428 97764 275434 97776
rect 282178 97764 282184 97776
rect 275428 97736 282184 97764
rect 275428 97724 275434 97736
rect 282178 97724 282184 97736
rect 282236 97724 282242 97776
rect 282730 97724 282736 97776
rect 282788 97764 282794 97776
rect 359458 97764 359464 97776
rect 282788 97736 359464 97764
rect 282788 97724 282794 97736
rect 359458 97724 359464 97736
rect 359516 97724 359522 97776
rect 221182 97696 221188 97708
rect 209056 97668 210556 97696
rect 215266 97668 221188 97696
rect 119338 97588 119344 97640
rect 119396 97628 119402 97640
rect 210528 97628 210556 97668
rect 221182 97656 221188 97668
rect 221240 97656 221246 97708
rect 227714 97656 227720 97708
rect 227772 97696 227778 97708
rect 229554 97696 229560 97708
rect 227772 97668 229560 97696
rect 227772 97656 227778 97668
rect 229554 97656 229560 97668
rect 229612 97656 229618 97708
rect 247310 97656 247316 97708
rect 247368 97696 247374 97708
rect 253198 97696 253204 97708
rect 247368 97668 253204 97696
rect 247368 97656 247374 97668
rect 253198 97656 253204 97668
rect 253256 97656 253262 97708
rect 254026 97656 254032 97708
rect 254084 97696 254090 97708
rect 262766 97696 262772 97708
rect 254084 97668 262772 97696
rect 254084 97656 254090 97668
rect 262766 97656 262772 97668
rect 262824 97656 262830 97708
rect 262950 97656 262956 97708
rect 263008 97696 263014 97708
rect 267642 97696 267648 97708
rect 263008 97668 267648 97696
rect 263008 97656 263014 97668
rect 267642 97656 267648 97668
rect 267700 97656 267706 97708
rect 270586 97656 270592 97708
rect 270644 97696 270650 97708
rect 270644 97668 272932 97696
rect 270644 97656 270650 97668
rect 216766 97628 216772 97640
rect 119396 97600 210464 97628
rect 210528 97600 216772 97628
rect 119396 97588 119402 97600
rect 115198 97520 115204 97572
rect 115256 97560 115262 97572
rect 205726 97560 205732 97572
rect 115256 97532 205732 97560
rect 115256 97520 115262 97532
rect 205726 97520 205732 97532
rect 205784 97520 205790 97572
rect 210436 97560 210464 97600
rect 216766 97588 216772 97600
rect 216824 97588 216830 97640
rect 250438 97588 250444 97640
rect 250496 97628 250502 97640
rect 262858 97628 262864 97640
rect 250496 97600 262864 97628
rect 250496 97588 250502 97600
rect 262858 97588 262864 97600
rect 262916 97588 262922 97640
rect 265802 97588 265808 97640
rect 265860 97628 265866 97640
rect 272702 97628 272708 97640
rect 265860 97600 272708 97628
rect 265860 97588 265866 97600
rect 272702 97588 272708 97600
rect 272760 97588 272766 97640
rect 272904 97628 272932 97668
rect 272978 97656 272984 97708
rect 273036 97696 273042 97708
rect 273036 97668 282224 97696
rect 273036 97656 273042 97668
rect 277302 97628 277308 97640
rect 272904 97600 277308 97628
rect 277302 97588 277308 97600
rect 277360 97588 277366 97640
rect 277762 97588 277768 97640
rect 277820 97628 277826 97640
rect 281994 97628 282000 97640
rect 277820 97600 282000 97628
rect 277820 97588 277826 97600
rect 281994 97588 282000 97600
rect 282052 97588 282058 97640
rect 282196 97628 282224 97668
rect 282270 97656 282276 97708
rect 282328 97696 282334 97708
rect 363598 97696 363604 97708
rect 282328 97668 363604 97696
rect 282328 97656 282334 97668
rect 363598 97656 363604 97668
rect 363656 97656 363662 97708
rect 370498 97628 370504 97640
rect 282196 97600 370504 97628
rect 370498 97588 370504 97600
rect 370556 97588 370562 97640
rect 218606 97560 218612 97572
rect 210436 97532 218612 97560
rect 218606 97520 218612 97532
rect 218664 97520 218670 97572
rect 218790 97520 218796 97572
rect 218848 97560 218854 97572
rect 224954 97560 224960 97572
rect 218848 97532 224960 97560
rect 218848 97520 218854 97532
rect 224954 97520 224960 97532
rect 225012 97520 225018 97572
rect 247494 97520 247500 97572
rect 247552 97560 247558 97572
rect 258718 97560 258724 97572
rect 247552 97532 258724 97560
rect 247552 97520 247558 97532
rect 258718 97520 258724 97532
rect 258776 97520 258782 97572
rect 262582 97520 262588 97572
rect 262640 97560 262646 97572
rect 369118 97560 369124 97572
rect 262640 97532 369124 97560
rect 262640 97520 262646 97532
rect 369118 97520 369124 97532
rect 369176 97520 369182 97572
rect 200206 97452 200212 97504
rect 200264 97492 200270 97504
rect 200942 97492 200948 97504
rect 200264 97464 200948 97492
rect 200264 97452 200270 97464
rect 200942 97452 200948 97464
rect 201000 97452 201006 97504
rect 203334 97452 203340 97504
rect 203392 97492 203398 97504
rect 206646 97492 206652 97504
rect 203392 97464 206652 97492
rect 203392 97452 203398 97464
rect 206646 97452 206652 97464
rect 206704 97452 206710 97504
rect 212534 97452 212540 97504
rect 212592 97492 212598 97504
rect 224218 97492 224224 97504
rect 212592 97464 224224 97492
rect 212592 97452 212598 97464
rect 224218 97452 224224 97464
rect 224276 97452 224282 97504
rect 257430 97452 257436 97504
rect 257488 97492 257494 97504
rect 263042 97492 263048 97504
rect 257488 97464 263048 97492
rect 257488 97452 257494 97464
rect 263042 97452 263048 97464
rect 263100 97452 263106 97504
rect 267734 97452 267740 97504
rect 267792 97492 267798 97504
rect 273254 97492 273260 97504
rect 267792 97464 273260 97492
rect 267792 97452 267798 97464
rect 273254 97452 273260 97464
rect 273312 97452 273318 97504
rect 278958 97452 278964 97504
rect 279016 97492 279022 97504
rect 281994 97492 282000 97504
rect 279016 97464 282000 97492
rect 279016 97452 279022 97464
rect 281994 97452 282000 97464
rect 282052 97452 282058 97504
rect 282178 97452 282184 97504
rect 282236 97492 282242 97504
rect 425698 97492 425704 97504
rect 282236 97464 425704 97492
rect 282236 97452 282242 97464
rect 425698 97452 425704 97464
rect 425756 97452 425762 97504
rect 97258 97384 97264 97436
rect 97316 97424 97322 97436
rect 215570 97424 215576 97436
rect 97316 97396 206692 97424
rect 97316 97384 97322 97396
rect 58618 97316 58624 97368
rect 58676 97356 58682 97368
rect 206002 97356 206008 97368
rect 58676 97328 206008 97356
rect 58676 97316 58682 97328
rect 206002 97316 206008 97328
rect 206060 97316 206066 97368
rect 206664 97356 206692 97396
rect 207032 97396 215576 97424
rect 207032 97356 207060 97396
rect 215570 97384 215576 97396
rect 215628 97384 215634 97436
rect 218054 97384 218060 97436
rect 218112 97424 218118 97436
rect 232498 97424 232504 97436
rect 218112 97396 232504 97424
rect 218112 97384 218118 97396
rect 232498 97384 232504 97396
rect 232556 97384 232562 97436
rect 244458 97384 244464 97436
rect 244516 97424 244522 97436
rect 248414 97424 248420 97436
rect 244516 97396 248420 97424
rect 244516 97384 244522 97396
rect 248414 97384 248420 97396
rect 248472 97384 248478 97436
rect 256970 97424 256976 97436
rect 252664 97396 256976 97424
rect 206664 97328 207060 97356
rect 208118 97316 208124 97368
rect 208176 97356 208182 97368
rect 227806 97356 227812 97368
rect 208176 97328 227812 97356
rect 208176 97316 208182 97328
rect 227806 97316 227812 97328
rect 227864 97316 227870 97368
rect 243262 97316 243268 97368
rect 243320 97356 243326 97368
rect 252664 97356 252692 97396
rect 256970 97384 256976 97396
rect 257028 97384 257034 97436
rect 263410 97384 263416 97436
rect 263468 97424 263474 97436
rect 271322 97424 271328 97436
rect 263468 97396 271328 97424
rect 263468 97384 263474 97396
rect 271322 97384 271328 97396
rect 271380 97384 271386 97436
rect 276566 97384 276572 97436
rect 276624 97424 276630 97436
rect 429838 97424 429844 97436
rect 276624 97396 429844 97424
rect 276624 97384 276630 97396
rect 429838 97384 429844 97396
rect 429896 97384 429902 97436
rect 243320 97328 252692 97356
rect 243320 97316 243326 97328
rect 253290 97316 253296 97368
rect 253348 97356 253354 97368
rect 258350 97356 258356 97368
rect 253348 97328 258356 97356
rect 253348 97316 253354 97328
rect 258350 97316 258356 97328
rect 258408 97316 258414 97368
rect 260466 97316 260472 97368
rect 260524 97356 260530 97368
rect 276658 97356 276664 97368
rect 260524 97328 276664 97356
rect 260524 97316 260530 97328
rect 276658 97316 276664 97328
rect 276716 97316 276722 97368
rect 276750 97316 276756 97368
rect 276808 97356 276814 97368
rect 277118 97356 277124 97368
rect 276808 97328 277124 97356
rect 276808 97316 276814 97328
rect 277118 97316 277124 97328
rect 277176 97316 277182 97368
rect 282270 97356 282276 97368
rect 277366 97328 282276 97356
rect 39942 97248 39948 97300
rect 40000 97288 40006 97300
rect 203334 97288 203340 97300
rect 40000 97260 203340 97288
rect 40000 97248 40006 97260
rect 203334 97248 203340 97260
rect 203392 97248 203398 97300
rect 206922 97248 206928 97300
rect 206980 97288 206986 97300
rect 227162 97288 227168 97300
rect 206980 97260 227168 97288
rect 206980 97248 206986 97260
rect 227162 97248 227168 97260
rect 227220 97248 227226 97300
rect 227622 97248 227628 97300
rect 227680 97288 227686 97300
rect 238294 97288 238300 97300
rect 227680 97260 238300 97288
rect 227680 97248 227686 97260
rect 238294 97248 238300 97260
rect 238352 97248 238358 97300
rect 246298 97248 246304 97300
rect 246356 97288 246362 97300
rect 271046 97288 271052 97300
rect 246356 97260 271052 97288
rect 246356 97248 246362 97260
rect 271046 97248 271052 97260
rect 271104 97248 271110 97300
rect 272426 97248 272432 97300
rect 272484 97288 272490 97300
rect 277366 97288 277394 97328
rect 282270 97316 282276 97328
rect 282328 97316 282334 97368
rect 285048 97328 285720 97356
rect 272484 97260 277394 97288
rect 272484 97248 272490 97260
rect 281074 97248 281080 97300
rect 281132 97288 281138 97300
rect 281350 97288 281356 97300
rect 281132 97260 281356 97288
rect 281132 97248 281138 97260
rect 281350 97248 281356 97260
rect 281408 97248 281414 97300
rect 281994 97248 282000 97300
rect 282052 97288 282058 97300
rect 285048 97288 285076 97328
rect 282052 97260 285076 97288
rect 282052 97248 282058 97260
rect 285122 97248 285128 97300
rect 285180 97288 285186 97300
rect 285582 97288 285588 97300
rect 285180 97260 285588 97288
rect 285180 97248 285186 97260
rect 285582 97248 285588 97260
rect 285640 97248 285646 97300
rect 285692 97288 285720 97328
rect 285858 97316 285864 97368
rect 285916 97356 285922 97368
rect 436738 97356 436744 97368
rect 285916 97328 436744 97356
rect 285916 97316 285922 97328
rect 436738 97316 436744 97328
rect 436796 97316 436802 97368
rect 443638 97288 443644 97300
rect 285692 97260 443644 97288
rect 443638 97248 443644 97260
rect 443696 97248 443702 97300
rect 142798 97180 142804 97232
rect 142856 97220 142862 97232
rect 208854 97220 208860 97232
rect 142856 97192 208860 97220
rect 142856 97180 142862 97192
rect 208854 97180 208860 97192
rect 208912 97180 208918 97232
rect 208946 97180 208952 97232
rect 209004 97220 209010 97232
rect 220998 97220 221004 97232
rect 209004 97192 221004 97220
rect 209004 97180 209010 97192
rect 220998 97180 221004 97192
rect 221056 97180 221062 97232
rect 248414 97180 248420 97232
rect 248472 97220 248478 97232
rect 260098 97220 260104 97232
rect 248472 97192 260104 97220
rect 248472 97180 248478 97192
rect 260098 97180 260104 97192
rect 260156 97180 260162 97232
rect 267274 97180 267280 97232
rect 267332 97220 267338 97232
rect 267332 97192 267734 97220
rect 267332 97180 267338 97192
rect 196618 97112 196624 97164
rect 196676 97152 196682 97164
rect 217962 97152 217968 97164
rect 196676 97124 217968 97152
rect 196676 97112 196682 97124
rect 217962 97112 217968 97124
rect 218020 97112 218026 97164
rect 219710 97112 219716 97164
rect 219768 97152 219774 97164
rect 220354 97152 220360 97164
rect 219768 97124 220360 97152
rect 219768 97112 219774 97124
rect 220354 97112 220360 97124
rect 220412 97112 220418 97164
rect 231854 97112 231860 97164
rect 231912 97152 231918 97164
rect 237742 97152 237748 97164
rect 231912 97124 237748 97152
rect 231912 97112 231918 97124
rect 237742 97112 237748 97124
rect 237800 97112 237806 97164
rect 240042 97112 240048 97164
rect 240100 97152 240106 97164
rect 242710 97152 242716 97164
rect 240100 97124 242716 97152
rect 240100 97112 240106 97124
rect 242710 97112 242716 97124
rect 242768 97112 242774 97164
rect 261018 97112 261024 97164
rect 261076 97152 261082 97164
rect 267706 97152 267734 97192
rect 268838 97180 268844 97232
rect 268896 97220 268902 97232
rect 269022 97220 269028 97232
rect 268896 97192 269028 97220
rect 268896 97180 268902 97192
rect 269022 97180 269028 97192
rect 269080 97180 269086 97232
rect 270034 97180 270040 97232
rect 270092 97220 270098 97232
rect 271138 97220 271144 97232
rect 270092 97192 271144 97220
rect 270092 97180 270098 97192
rect 271138 97180 271144 97192
rect 271196 97180 271202 97232
rect 274174 97180 274180 97232
rect 274232 97220 274238 97232
rect 274542 97220 274548 97232
rect 274232 97192 274548 97220
rect 274232 97180 274238 97192
rect 274542 97180 274548 97192
rect 274600 97180 274606 97232
rect 275554 97180 275560 97232
rect 275612 97220 275618 97232
rect 275922 97220 275928 97232
rect 275612 97192 275928 97220
rect 275612 97180 275618 97192
rect 275922 97180 275928 97192
rect 275980 97180 275986 97232
rect 276014 97180 276020 97232
rect 276072 97220 276078 97232
rect 323578 97220 323584 97232
rect 276072 97192 323584 97220
rect 276072 97180 276078 97192
rect 323578 97180 323584 97192
rect 323636 97180 323642 97232
rect 298002 97152 298008 97164
rect 261076 97124 266860 97152
rect 267706 97124 298008 97152
rect 261076 97112 261082 97124
rect 192478 97044 192484 97096
rect 192536 97084 192542 97096
rect 202690 97084 202696 97096
rect 192536 97056 202696 97084
rect 192536 97044 192542 97056
rect 202690 97044 202696 97056
rect 202748 97044 202754 97096
rect 202782 97044 202788 97096
rect 202840 97084 202846 97096
rect 205450 97084 205456 97096
rect 202840 97056 205456 97084
rect 202840 97044 202846 97056
rect 205450 97044 205456 97056
rect 205508 97044 205514 97096
rect 205726 97044 205732 97096
rect 205784 97084 205790 97096
rect 219158 97084 219164 97096
rect 205784 97056 219164 97084
rect 205784 97044 205790 97056
rect 219158 97044 219164 97056
rect 219216 97044 219222 97096
rect 241330 97044 241336 97096
rect 241388 97084 241394 97096
rect 242158 97084 242164 97096
rect 241388 97056 242164 97084
rect 241388 97044 241394 97056
rect 242158 97044 242164 97056
rect 242216 97044 242222 97096
rect 246666 97044 246672 97096
rect 246724 97084 246730 97096
rect 246850 97084 246856 97096
rect 246724 97056 246856 97084
rect 246724 97044 246730 97056
rect 246850 97044 246856 97056
rect 246908 97044 246914 97096
rect 253474 97044 253480 97096
rect 253532 97084 253538 97096
rect 253750 97084 253756 97096
rect 253532 97056 253756 97084
rect 253532 97044 253538 97056
rect 253750 97044 253756 97056
rect 253808 97044 253814 97096
rect 255038 97044 255044 97096
rect 255096 97084 255102 97096
rect 255096 97056 255268 97084
rect 255096 97044 255102 97056
rect 197998 96976 198004 97028
rect 198056 97016 198062 97028
rect 211430 97016 211436 97028
rect 198056 96988 202736 97016
rect 198056 96976 198062 96988
rect 195238 96908 195244 96960
rect 195296 96948 195302 96960
rect 201862 96948 201868 96960
rect 195296 96920 201868 96948
rect 195296 96908 195302 96920
rect 201862 96908 201868 96920
rect 201920 96908 201926 96960
rect 201954 96908 201960 96960
rect 202012 96948 202018 96960
rect 202506 96948 202512 96960
rect 202012 96920 202512 96948
rect 202012 96908 202018 96920
rect 202506 96908 202512 96920
rect 202564 96908 202570 96960
rect 202708 96948 202736 96988
rect 202984 96988 211436 97016
rect 202984 96948 203012 96988
rect 211430 96976 211436 96988
rect 211488 96976 211494 97028
rect 241698 96976 241704 97028
rect 241756 97016 241762 97028
rect 242526 97016 242532 97028
rect 241756 96988 242532 97016
rect 241756 96976 241762 96988
rect 242526 96976 242532 96988
rect 242584 96976 242590 97028
rect 250070 96976 250076 97028
rect 250128 97016 250134 97028
rect 250714 97016 250720 97028
rect 250128 96988 250720 97016
rect 250128 96976 250134 96988
rect 250714 96976 250720 96988
rect 250772 96976 250778 97028
rect 251266 96976 251272 97028
rect 251324 97016 251330 97028
rect 252186 97016 252192 97028
rect 251324 96988 252192 97016
rect 251324 96976 251330 96988
rect 252186 96976 252192 96988
rect 252244 96976 252250 97028
rect 252278 96976 252284 97028
rect 252336 97016 252342 97028
rect 252462 97016 252468 97028
rect 252336 96988 252468 97016
rect 252336 96976 252342 96988
rect 252462 96976 252468 96988
rect 252520 96976 252526 97028
rect 254670 96976 254676 97028
rect 254728 97016 254734 97028
rect 255130 97016 255136 97028
rect 254728 96988 255136 97016
rect 254728 96976 254734 96988
rect 255130 96976 255136 96988
rect 255188 96976 255194 97028
rect 202708 96920 203012 96948
rect 208854 96908 208860 96960
rect 208912 96948 208918 96960
rect 212626 96948 212632 96960
rect 208912 96920 212632 96948
rect 208912 96908 208918 96920
rect 212626 96908 212632 96920
rect 212684 96908 212690 96960
rect 215754 96908 215760 96960
rect 215812 96948 215818 96960
rect 216306 96948 216312 96960
rect 215812 96920 216312 96948
rect 215812 96908 215818 96920
rect 216306 96908 216312 96920
rect 216364 96908 216370 96960
rect 216858 96908 216864 96960
rect 216916 96948 216922 96960
rect 217134 96948 217140 96960
rect 216916 96920 217140 96948
rect 216916 96908 216922 96920
rect 217134 96908 217140 96920
rect 217192 96908 217198 96960
rect 219710 96908 219716 96960
rect 219768 96948 219774 96960
rect 220446 96948 220452 96960
rect 219768 96920 220452 96948
rect 219768 96908 219774 96920
rect 220446 96908 220452 96920
rect 220504 96908 220510 96960
rect 221458 96908 221464 96960
rect 221516 96948 221522 96960
rect 221918 96948 221924 96960
rect 221516 96920 221924 96948
rect 221516 96908 221522 96920
rect 221918 96908 221924 96920
rect 221976 96908 221982 96960
rect 222286 96908 222292 96960
rect 222344 96948 222350 96960
rect 222930 96948 222936 96960
rect 222344 96920 222936 96948
rect 222344 96908 222350 96920
rect 222930 96908 222936 96920
rect 222988 96908 222994 96960
rect 234706 96908 234712 96960
rect 234764 96948 234770 96960
rect 235442 96948 235448 96960
rect 234764 96920 235448 96948
rect 234764 96908 234770 96920
rect 235442 96908 235448 96920
rect 235500 96908 235506 96960
rect 236454 96908 236460 96960
rect 236512 96948 236518 96960
rect 237190 96948 237196 96960
rect 236512 96920 237196 96948
rect 236512 96908 236518 96920
rect 237190 96908 237196 96920
rect 237248 96908 237254 96960
rect 237650 96908 237656 96960
rect 237708 96948 237714 96960
rect 238386 96948 238392 96960
rect 237708 96920 238392 96948
rect 237708 96908 237714 96920
rect 238386 96908 238392 96920
rect 238444 96908 238450 96960
rect 239030 96908 239036 96960
rect 239088 96948 239094 96960
rect 239398 96948 239404 96960
rect 239088 96920 239404 96948
rect 239088 96908 239094 96920
rect 239398 96908 239404 96920
rect 239456 96908 239462 96960
rect 240318 96908 240324 96960
rect 240376 96948 240382 96960
rect 240778 96948 240784 96960
rect 240376 96920 240784 96948
rect 240376 96908 240382 96920
rect 240778 96908 240784 96920
rect 240836 96908 240842 96960
rect 241514 96908 241520 96960
rect 241572 96948 241578 96960
rect 242434 96948 242440 96960
rect 241572 96920 242440 96948
rect 241572 96908 241578 96920
rect 242434 96908 242440 96920
rect 242492 96908 242498 96960
rect 243722 96908 243728 96960
rect 243780 96948 243786 96960
rect 244090 96948 244096 96960
rect 243780 96920 244096 96948
rect 243780 96908 243786 96920
rect 244090 96908 244096 96920
rect 244148 96908 244154 96960
rect 244734 96908 244740 96960
rect 244792 96948 244798 96960
rect 245378 96948 245384 96960
rect 244792 96920 245384 96948
rect 244792 96908 244798 96920
rect 245378 96908 245384 96920
rect 245436 96908 245442 96960
rect 245930 96908 245936 96960
rect 245988 96948 245994 96960
rect 246574 96948 246580 96960
rect 245988 96920 246580 96948
rect 245988 96908 245994 96920
rect 246574 96908 246580 96920
rect 246632 96908 246638 96960
rect 247126 96908 247132 96960
rect 247184 96948 247190 96960
rect 248230 96948 248236 96960
rect 247184 96920 248236 96948
rect 247184 96908 247190 96920
rect 248230 96908 248236 96920
rect 248288 96908 248294 96960
rect 248506 96908 248512 96960
rect 248564 96948 248570 96960
rect 249334 96948 249340 96960
rect 248564 96920 249340 96948
rect 248564 96908 248570 96920
rect 249334 96908 249340 96920
rect 249392 96908 249398 96960
rect 250622 96908 250628 96960
rect 250680 96948 250686 96960
rect 250990 96948 250996 96960
rect 250680 96920 250996 96948
rect 250680 96908 250686 96920
rect 250990 96908 250996 96920
rect 251048 96908 251054 96960
rect 251450 96908 251456 96960
rect 251508 96948 251514 96960
rect 252002 96948 252008 96960
rect 251508 96920 252008 96948
rect 251508 96908 251514 96920
rect 252002 96908 252008 96920
rect 252060 96908 252066 96960
rect 252646 96908 252652 96960
rect 252704 96948 252710 96960
rect 253658 96948 253664 96960
rect 252704 96920 253664 96948
rect 252704 96908 252710 96920
rect 253658 96908 253664 96920
rect 253716 96908 253722 96960
rect 254210 96908 254216 96960
rect 254268 96948 254274 96960
rect 255038 96948 255044 96960
rect 254268 96920 255044 96948
rect 254268 96908 254274 96920
rect 255038 96908 255044 96920
rect 255096 96908 255102 96960
rect 199378 96840 199384 96892
rect 199436 96880 199442 96892
rect 202782 96880 202788 96892
rect 199436 96852 202788 96880
rect 199436 96840 199442 96852
rect 202782 96840 202788 96852
rect 202840 96840 202846 96892
rect 203518 96840 203524 96892
rect 203576 96880 203582 96892
rect 207198 96880 207204 96892
rect 203576 96852 207204 96880
rect 203576 96840 203582 96852
rect 207198 96840 207204 96852
rect 207256 96840 207262 96892
rect 222470 96840 222476 96892
rect 222528 96880 222534 96892
rect 223298 96880 223304 96892
rect 222528 96852 223304 96880
rect 222528 96840 222534 96852
rect 223298 96840 223304 96852
rect 223356 96840 223362 96892
rect 234614 96840 234620 96892
rect 234672 96880 234678 96892
rect 235810 96880 235816 96892
rect 234672 96852 235816 96880
rect 234672 96840 234678 96852
rect 235810 96840 235816 96852
rect 235868 96840 235874 96892
rect 240226 96840 240232 96892
rect 240284 96880 240290 96892
rect 240962 96880 240968 96892
rect 240284 96852 240968 96880
rect 240284 96840 240290 96852
rect 240962 96840 240968 96852
rect 241020 96840 241026 96892
rect 242342 96840 242348 96892
rect 242400 96880 242406 96892
rect 242802 96880 242808 96892
rect 242400 96852 242808 96880
rect 242400 96840 242406 96852
rect 242802 96840 242808 96852
rect 242860 96840 242866 96892
rect 245102 96840 245108 96892
rect 245160 96880 245166 96892
rect 245470 96880 245476 96892
rect 245160 96852 245476 96880
rect 245160 96840 245166 96852
rect 245470 96840 245476 96852
rect 245528 96840 245534 96892
rect 246114 96840 246120 96892
rect 246172 96880 246178 96892
rect 246942 96880 246948 96892
rect 246172 96852 246948 96880
rect 246172 96840 246178 96852
rect 246942 96840 246948 96852
rect 247000 96840 247006 96892
rect 248690 96840 248696 96892
rect 248748 96880 248754 96892
rect 249518 96880 249524 96892
rect 248748 96852 249524 96880
rect 248748 96840 248754 96852
rect 249518 96840 249524 96852
rect 249576 96840 249582 96892
rect 250254 96840 250260 96892
rect 250312 96880 250318 96892
rect 250806 96880 250812 96892
rect 250312 96852 250812 96880
rect 250312 96840 250318 96852
rect 250806 96840 250812 96852
rect 250864 96840 250870 96892
rect 251818 96840 251824 96892
rect 251876 96880 251882 96892
rect 252278 96880 252284 96892
rect 251876 96852 252284 96880
rect 251876 96840 251882 96852
rect 252278 96840 252284 96852
rect 252336 96840 252342 96892
rect 255240 96880 255268 97056
rect 265894 97044 265900 97096
rect 265952 97084 265958 97096
rect 266170 97084 266176 97096
rect 265952 97056 266176 97084
rect 265952 97044 265958 97056
rect 266170 97044 266176 97056
rect 266228 97044 266234 97096
rect 266832 97084 266860 97124
rect 298002 97112 298008 97124
rect 298060 97112 298066 97164
rect 302878 97152 302884 97164
rect 302206 97124 302884 97152
rect 266832 97056 267136 97084
rect 256050 96976 256056 97028
rect 256108 97016 256114 97028
rect 256418 97016 256424 97028
rect 256108 96988 256424 97016
rect 256108 96976 256114 96988
rect 256418 96976 256424 96988
rect 256476 96976 256482 97028
rect 257246 96976 257252 97028
rect 257304 97016 257310 97028
rect 257890 97016 257896 97028
rect 257304 96988 257896 97016
rect 257304 96976 257310 96988
rect 257890 96976 257896 96988
rect 257948 96976 257954 97028
rect 258074 96976 258080 97028
rect 258132 97016 258138 97028
rect 259086 97016 259092 97028
rect 258132 96988 259092 97016
rect 258132 96976 258138 96988
rect 259086 96976 259092 96988
rect 259144 96976 259150 97028
rect 261754 96976 261760 97028
rect 261812 97016 261818 97028
rect 262030 97016 262036 97028
rect 261812 96988 262036 97016
rect 261812 96976 261818 96988
rect 262030 96976 262036 96988
rect 262088 96976 262094 97028
rect 263594 96976 263600 97028
rect 263652 97016 263658 97028
rect 264790 97016 264796 97028
rect 263652 96988 264796 97016
rect 263652 96976 263658 96988
rect 264790 96976 264796 96988
rect 264848 96976 264854 97028
rect 265434 96976 265440 97028
rect 265492 97016 265498 97028
rect 266998 97016 267004 97028
rect 265492 96988 267004 97016
rect 265492 96976 265498 96988
rect 266998 96976 267004 96988
rect 267056 96976 267062 97028
rect 267108 97016 267136 97056
rect 267182 97044 267188 97096
rect 267240 97084 267246 97096
rect 267550 97084 267556 97096
rect 267240 97056 267556 97084
rect 267240 97044 267246 97056
rect 267550 97044 267556 97056
rect 267608 97044 267614 97096
rect 267642 97044 267648 97096
rect 267700 97084 267706 97096
rect 302206 97084 302234 97124
rect 302878 97112 302884 97124
rect 302936 97112 302942 97164
rect 267700 97056 302234 97084
rect 267700 97044 267706 97056
rect 300118 97016 300124 97028
rect 267108 96988 300124 97016
rect 300118 96976 300124 96988
rect 300176 96976 300182 97028
rect 255682 96908 255688 96960
rect 255740 96948 255746 96960
rect 256142 96948 256148 96960
rect 255740 96920 256148 96948
rect 255740 96908 255746 96920
rect 256142 96908 256148 96920
rect 256200 96908 256206 96960
rect 256326 96908 256332 96960
rect 256384 96948 256390 96960
rect 256602 96948 256608 96960
rect 256384 96920 256608 96948
rect 256384 96908 256390 96920
rect 256602 96908 256608 96920
rect 256660 96908 256666 96960
rect 257614 96908 257620 96960
rect 257672 96948 257678 96960
rect 257982 96948 257988 96960
rect 257672 96920 257988 96948
rect 257672 96908 257678 96920
rect 257982 96908 257988 96920
rect 258040 96908 258046 96960
rect 258442 96908 258448 96960
rect 258500 96948 258506 96960
rect 258994 96948 259000 96960
rect 258500 96920 259000 96948
rect 258500 96908 258506 96920
rect 258994 96908 259000 96920
rect 259052 96908 259058 96960
rect 259454 96908 259460 96960
rect 259512 96948 259518 96960
rect 260282 96948 260288 96960
rect 259512 96920 260288 96948
rect 259512 96908 259518 96920
rect 260282 96908 260288 96920
rect 260340 96908 260346 96960
rect 261202 96908 261208 96960
rect 261260 96948 261266 96960
rect 261846 96948 261852 96960
rect 261260 96920 261852 96948
rect 261260 96908 261266 96920
rect 261846 96908 261852 96920
rect 261904 96908 261910 96960
rect 264054 96908 264060 96960
rect 264112 96948 264118 96960
rect 264514 96948 264520 96960
rect 264112 96920 264520 96948
rect 264112 96908 264118 96920
rect 264514 96908 264520 96920
rect 264572 96908 264578 96960
rect 265250 96908 265256 96960
rect 265308 96948 265314 96960
rect 265986 96948 265992 96960
rect 265308 96920 265992 96948
rect 265308 96908 265314 96920
rect 265986 96908 265992 96920
rect 266044 96908 266050 96960
rect 266814 96908 266820 96960
rect 266872 96948 266878 96960
rect 267366 96948 267372 96960
rect 266872 96920 267372 96948
rect 266872 96908 266878 96920
rect 267366 96908 267372 96920
rect 267424 96908 267430 96960
rect 268010 96908 268016 96960
rect 268068 96948 268074 96960
rect 268654 96948 268660 96960
rect 268068 96920 268660 96948
rect 268068 96908 268074 96920
rect 268654 96908 268660 96920
rect 268712 96908 268718 96960
rect 269758 96908 269764 96960
rect 269816 96948 269822 96960
rect 270218 96948 270224 96960
rect 269816 96920 270224 96948
rect 269816 96908 269822 96920
rect 270218 96908 270224 96920
rect 270276 96908 270282 96960
rect 271230 96908 271236 96960
rect 271288 96948 271294 96960
rect 271782 96948 271788 96960
rect 271288 96920 271788 96948
rect 271288 96908 271294 96920
rect 271782 96908 271788 96920
rect 271840 96908 271846 96960
rect 272610 96908 272616 96960
rect 272668 96948 272674 96960
rect 272886 96948 272892 96960
rect 272668 96920 272892 96948
rect 272668 96908 272674 96920
rect 272886 96908 272892 96920
rect 272944 96908 272950 96960
rect 273254 96908 273260 96960
rect 273312 96948 273318 96960
rect 298830 96948 298836 96960
rect 273312 96920 298836 96948
rect 273312 96908 273318 96920
rect 298830 96908 298836 96920
rect 298888 96908 298894 96960
rect 255240 96852 255360 96880
rect 98638 96772 98644 96824
rect 98696 96812 98702 96824
rect 204070 96812 204076 96824
rect 98696 96784 200114 96812
rect 98696 96772 98702 96784
rect 200086 96676 200114 96784
rect 200316 96784 204076 96812
rect 200316 96676 200344 96784
rect 204070 96772 204076 96784
rect 204128 96772 204134 96824
rect 215478 96772 215484 96824
rect 215536 96812 215542 96824
rect 216490 96812 216496 96824
rect 215536 96784 216496 96812
rect 215536 96772 215542 96784
rect 216490 96772 216496 96784
rect 216548 96772 216554 96824
rect 217134 96772 217140 96824
rect 217192 96812 217198 96824
rect 217686 96812 217692 96824
rect 217192 96784 217692 96812
rect 217192 96772 217198 96784
rect 217686 96772 217692 96784
rect 217744 96772 217750 96824
rect 218238 96772 218244 96824
rect 218296 96812 218302 96824
rect 218882 96812 218888 96824
rect 218296 96784 218888 96812
rect 218296 96772 218302 96784
rect 218882 96772 218888 96784
rect 218940 96772 218946 96824
rect 219434 96772 219440 96824
rect 219492 96812 219498 96824
rect 220446 96812 220452 96824
rect 219492 96784 220452 96812
rect 219492 96772 219498 96784
rect 220446 96772 220452 96784
rect 220504 96772 220510 96824
rect 221090 96772 221096 96824
rect 221148 96812 221154 96824
rect 221642 96812 221648 96824
rect 221148 96784 221648 96812
rect 221148 96772 221154 96784
rect 221642 96772 221648 96784
rect 221700 96772 221706 96824
rect 222286 96772 222292 96824
rect 222344 96812 222350 96824
rect 223114 96812 223120 96824
rect 222344 96784 223120 96812
rect 222344 96772 222350 96784
rect 223114 96772 223120 96784
rect 223172 96772 223178 96824
rect 231578 96772 231584 96824
rect 231636 96812 231642 96824
rect 237098 96812 237104 96824
rect 231636 96784 237104 96812
rect 231636 96772 231642 96784
rect 237098 96772 237104 96784
rect 237156 96772 237162 96824
rect 240686 96772 240692 96824
rect 240744 96812 240750 96824
rect 241330 96812 241336 96824
rect 240744 96784 241336 96812
rect 240744 96772 240750 96784
rect 241330 96772 241336 96784
rect 241388 96772 241394 96824
rect 241882 96772 241888 96824
rect 241940 96812 241946 96824
rect 242710 96812 242716 96824
rect 241940 96784 242716 96812
rect 241940 96772 241946 96784
rect 242710 96772 242716 96784
rect 242768 96772 242774 96824
rect 245654 96772 245660 96824
rect 245712 96812 245718 96824
rect 246758 96812 246764 96824
rect 245712 96784 246764 96812
rect 245712 96772 245718 96784
rect 246758 96772 246764 96784
rect 246816 96772 246822 96824
rect 253382 96772 253388 96824
rect 253440 96812 253446 96824
rect 253842 96812 253848 96824
rect 253440 96784 253848 96812
rect 253440 96772 253446 96784
rect 253842 96772 253848 96784
rect 253900 96772 253906 96824
rect 254762 96772 254768 96824
rect 254820 96812 254826 96824
rect 255222 96812 255228 96824
rect 254820 96784 255228 96812
rect 254820 96772 254826 96784
rect 255222 96772 255228 96784
rect 255280 96772 255286 96824
rect 201862 96704 201868 96756
rect 201920 96744 201926 96756
rect 206462 96744 206468 96756
rect 201920 96716 206468 96744
rect 201920 96704 201926 96716
rect 206462 96704 206468 96716
rect 206520 96704 206526 96756
rect 244274 96704 244280 96756
rect 244332 96744 244338 96756
rect 245470 96744 245476 96756
rect 244332 96716 245476 96744
rect 244332 96704 244338 96716
rect 245470 96704 245476 96716
rect 245528 96704 245534 96756
rect 200086 96648 200344 96676
rect 202690 96636 202696 96688
rect 202748 96676 202754 96688
rect 208394 96676 208400 96688
rect 202748 96648 208400 96676
rect 202748 96636 202754 96648
rect 208394 96636 208400 96648
rect 208452 96636 208458 96688
rect 210418 96636 210424 96688
rect 210476 96676 210482 96688
rect 216214 96676 216220 96688
rect 210476 96648 216220 96676
rect 210476 96636 210482 96648
rect 216214 96636 216220 96648
rect 216272 96636 216278 96688
rect 243078 96636 243084 96688
rect 243136 96676 243142 96688
rect 246298 96676 246304 96688
rect 243136 96648 246304 96676
rect 243136 96636 243142 96648
rect 246298 96636 246304 96648
rect 246356 96636 246362 96688
rect 186958 96568 186964 96620
rect 187016 96608 187022 96620
rect 231302 96608 231308 96620
rect 187016 96580 231308 96608
rect 187016 96568 187022 96580
rect 231302 96568 231308 96580
rect 231360 96568 231366 96620
rect 255332 96608 255360 96852
rect 257062 96840 257068 96892
rect 257120 96880 257126 96892
rect 257798 96880 257804 96892
rect 257120 96852 257804 96880
rect 257120 96840 257126 96852
rect 257798 96840 257804 96852
rect 257856 96840 257862 96892
rect 258810 96840 258816 96892
rect 258868 96880 258874 96892
rect 259362 96880 259368 96892
rect 258868 96852 259368 96880
rect 258868 96840 258874 96852
rect 259362 96840 259368 96852
rect 259420 96840 259426 96892
rect 259638 96840 259644 96892
rect 259696 96880 259702 96892
rect 260742 96880 260748 96892
rect 259696 96852 260748 96880
rect 259696 96840 259702 96852
rect 260742 96840 260748 96852
rect 260800 96840 260806 96892
rect 261662 96840 261668 96892
rect 261720 96880 261726 96892
rect 262950 96880 262956 96892
rect 261720 96852 262956 96880
rect 261720 96840 261726 96852
rect 262950 96840 262956 96852
rect 263008 96840 263014 96892
rect 264238 96840 264244 96892
rect 264296 96880 264302 96892
rect 264882 96880 264888 96892
rect 264296 96852 264888 96880
rect 264296 96840 264302 96852
rect 264882 96840 264888 96852
rect 264940 96840 264946 96892
rect 266630 96840 266636 96892
rect 266688 96880 266694 96892
rect 267642 96880 267648 96892
rect 266688 96852 267648 96880
rect 266688 96840 266694 96852
rect 267642 96840 267648 96852
rect 267700 96840 267706 96892
rect 267826 96840 267832 96892
rect 267884 96880 267890 96892
rect 268562 96880 268568 96892
rect 267884 96852 268568 96880
rect 267884 96840 267890 96852
rect 268562 96840 268568 96852
rect 268620 96840 268626 96892
rect 269574 96840 269580 96892
rect 269632 96880 269638 96892
rect 270310 96880 270316 96892
rect 269632 96852 270316 96880
rect 269632 96840 269638 96852
rect 270310 96840 270316 96852
rect 270368 96840 270374 96892
rect 271966 96840 271972 96892
rect 272024 96880 272030 96892
rect 273162 96880 273168 96892
rect 272024 96852 273168 96880
rect 272024 96840 272030 96852
rect 273162 96840 273168 96852
rect 273220 96840 273226 96892
rect 273272 96852 277256 96880
rect 255406 96772 255412 96824
rect 255464 96812 255470 96824
rect 256050 96812 256056 96824
rect 255464 96784 256056 96812
rect 255464 96772 255470 96784
rect 256050 96772 256056 96784
rect 256108 96772 256114 96824
rect 258258 96772 258264 96824
rect 258316 96812 258322 96824
rect 259178 96812 259184 96824
rect 258316 96784 259184 96812
rect 258316 96772 258322 96784
rect 259178 96772 259184 96784
rect 259236 96772 259242 96824
rect 260190 96772 260196 96824
rect 260248 96812 260254 96824
rect 260466 96812 260472 96824
rect 260248 96784 260472 96812
rect 260248 96772 260254 96784
rect 260466 96772 260472 96784
rect 260524 96772 260530 96824
rect 262398 96772 262404 96824
rect 262456 96812 262462 96824
rect 263318 96812 263324 96824
rect 262456 96784 263324 96812
rect 262456 96772 262462 96784
rect 263318 96772 263324 96784
rect 263376 96772 263382 96824
rect 263778 96772 263784 96824
rect 263836 96812 263842 96824
rect 264698 96812 264704 96824
rect 263836 96784 264704 96812
rect 263836 96772 263842 96784
rect 264698 96772 264704 96784
rect 264756 96772 264762 96824
rect 265618 96772 265624 96824
rect 265676 96812 265682 96824
rect 266170 96812 266176 96824
rect 265676 96784 266176 96812
rect 265676 96772 265682 96784
rect 266170 96772 266176 96784
rect 266228 96772 266234 96824
rect 266446 96772 266452 96824
rect 266504 96812 266510 96824
rect 267182 96812 267188 96824
rect 266504 96784 267188 96812
rect 266504 96772 266510 96784
rect 267182 96772 267188 96784
rect 267240 96772 267246 96824
rect 268378 96772 268384 96824
rect 268436 96812 268442 96824
rect 268930 96812 268936 96824
rect 268436 96784 268936 96812
rect 268436 96772 268442 96784
rect 268930 96772 268936 96784
rect 268988 96772 268994 96824
rect 269390 96772 269396 96824
rect 269448 96812 269454 96824
rect 270034 96812 270040 96824
rect 269448 96784 270040 96812
rect 269448 96772 269454 96784
rect 270034 96772 270040 96784
rect 270092 96772 270098 96824
rect 272150 96772 272156 96824
rect 272208 96812 272214 96824
rect 273070 96812 273076 96824
rect 272208 96784 273076 96812
rect 272208 96772 272214 96784
rect 273070 96772 273076 96784
rect 273128 96772 273134 96824
rect 260006 96704 260012 96756
rect 260064 96744 260070 96756
rect 260558 96744 260564 96756
rect 260064 96716 260564 96744
rect 260064 96704 260070 96716
rect 260558 96704 260564 96716
rect 260616 96704 260622 96756
rect 261386 96704 261392 96756
rect 261444 96744 261450 96756
rect 262030 96744 262036 96756
rect 261444 96716 262036 96744
rect 261444 96704 261450 96716
rect 262030 96704 262036 96716
rect 262088 96704 262094 96756
rect 262214 96704 262220 96756
rect 262272 96744 262278 96756
rect 263410 96744 263416 96756
rect 262272 96716 263416 96744
rect 262272 96704 262278 96716
rect 263410 96704 263416 96716
rect 263468 96704 263474 96756
rect 264974 96704 264980 96756
rect 265032 96744 265038 96756
rect 266078 96744 266084 96756
rect 265032 96716 266084 96744
rect 265032 96704 265038 96716
rect 266078 96704 266084 96716
rect 266136 96704 266142 96756
rect 269206 96704 269212 96756
rect 269264 96744 269270 96756
rect 270126 96744 270132 96756
rect 269264 96716 270132 96744
rect 269264 96704 269270 96716
rect 270126 96704 270132 96716
rect 270184 96704 270190 96756
rect 271874 96704 271880 96756
rect 271932 96744 271938 96756
rect 273272 96744 273300 96852
rect 274082 96772 274088 96824
rect 274140 96812 274146 96824
rect 274358 96812 274364 96824
rect 274140 96784 274364 96812
rect 274140 96772 274146 96784
rect 274358 96772 274364 96784
rect 274416 96772 274422 96824
rect 277228 96812 277256 96852
rect 277302 96840 277308 96892
rect 277360 96880 277366 96892
rect 278130 96880 278136 96892
rect 277360 96852 278136 96880
rect 277360 96840 277366 96852
rect 278130 96840 278136 96852
rect 278188 96840 278194 96892
rect 278314 96840 278320 96892
rect 278372 96880 278378 96892
rect 278498 96880 278504 96892
rect 278372 96852 278504 96880
rect 278372 96840 278378 96852
rect 278498 96840 278504 96852
rect 278556 96840 278562 96892
rect 279326 96840 279332 96892
rect 279384 96880 279390 96892
rect 279970 96880 279976 96892
rect 279384 96852 279976 96880
rect 279384 96840 279390 96852
rect 279970 96840 279976 96852
rect 280028 96840 280034 96892
rect 280522 96840 280528 96892
rect 280580 96880 280586 96892
rect 281166 96880 281172 96892
rect 280580 96852 281172 96880
rect 280580 96840 280586 96852
rect 281166 96840 281172 96852
rect 281224 96840 281230 96892
rect 281718 96840 281724 96892
rect 281776 96880 281782 96892
rect 282638 96880 282644 96892
rect 281776 96852 282644 96880
rect 281776 96840 281782 96852
rect 282638 96840 282644 96852
rect 282696 96840 282702 96892
rect 283742 96840 283748 96892
rect 283800 96880 283806 96892
rect 284110 96880 284116 96892
rect 283800 96852 284116 96880
rect 283800 96840 283806 96852
rect 284110 96840 284116 96852
rect 284168 96840 284174 96892
rect 284294 96840 284300 96892
rect 284352 96880 284358 96892
rect 285490 96880 285496 96892
rect 284352 96852 285496 96880
rect 284352 96840 284358 96852
rect 285490 96840 285496 96852
rect 285548 96840 285554 96892
rect 285950 96840 285956 96892
rect 286008 96880 286014 96892
rect 286686 96880 286692 96892
rect 286008 96852 286692 96880
rect 286008 96840 286014 96852
rect 286686 96840 286692 96852
rect 286744 96840 286750 96892
rect 307018 96880 307024 96892
rect 287026 96852 307024 96880
rect 277228 96784 277532 96812
rect 271932 96716 273300 96744
rect 271932 96704 271938 96716
rect 273346 96704 273352 96756
rect 273404 96744 273410 96756
rect 274634 96744 274640 96756
rect 273404 96716 274640 96744
rect 273404 96704 273410 96716
rect 274634 96704 274640 96716
rect 274692 96704 274698 96756
rect 275554 96704 275560 96756
rect 275612 96744 275618 96756
rect 275830 96744 275836 96756
rect 275612 96716 275836 96744
rect 275612 96704 275618 96716
rect 275830 96704 275836 96716
rect 275888 96704 275894 96756
rect 276198 96704 276204 96756
rect 276256 96744 276262 96756
rect 277302 96744 277308 96756
rect 276256 96716 277308 96744
rect 276256 96704 276262 96716
rect 277302 96704 277308 96716
rect 277360 96704 277366 96756
rect 260834 96636 260840 96688
rect 260892 96676 260898 96688
rect 261938 96676 261944 96688
rect 260892 96648 261944 96676
rect 260892 96636 260898 96648
rect 261938 96636 261944 96648
rect 261996 96636 262002 96688
rect 273622 96636 273628 96688
rect 273680 96676 273686 96688
rect 273680 96648 274404 96676
rect 273680 96636 273686 96648
rect 255332 96580 258074 96608
rect 161382 96500 161388 96552
rect 161440 96540 161446 96552
rect 206922 96540 206928 96552
rect 161440 96512 206928 96540
rect 161440 96500 161446 96512
rect 206922 96500 206928 96512
rect 206980 96500 206986 96552
rect 183462 96432 183468 96484
rect 183520 96472 183526 96484
rect 230750 96472 230756 96484
rect 183520 96444 230756 96472
rect 183520 96432 183526 96444
rect 230750 96432 230756 96444
rect 230808 96432 230814 96484
rect 258046 96472 258074 96580
rect 274376 96552 274404 96648
rect 274818 96636 274824 96688
rect 274876 96676 274882 96688
rect 274876 96648 275876 96676
rect 274876 96636 274882 96648
rect 275848 96552 275876 96648
rect 276382 96636 276388 96688
rect 276440 96676 276446 96688
rect 277210 96676 277216 96688
rect 276440 96648 277216 96676
rect 276440 96636 276446 96648
rect 277210 96636 277216 96648
rect 277268 96636 277274 96688
rect 277504 96676 277532 96784
rect 277946 96772 277952 96824
rect 278004 96812 278010 96824
rect 278682 96812 278688 96824
rect 278004 96784 278688 96812
rect 278004 96772 278010 96784
rect 278682 96772 278688 96784
rect 278740 96772 278746 96824
rect 278774 96772 278780 96824
rect 278832 96812 278838 96824
rect 279878 96812 279884 96824
rect 278832 96784 279884 96812
rect 278832 96772 278838 96784
rect 279878 96772 279884 96784
rect 279936 96772 279942 96824
rect 280338 96772 280344 96824
rect 280396 96812 280402 96824
rect 281258 96812 281264 96824
rect 280396 96784 281264 96812
rect 280396 96772 280402 96784
rect 281258 96772 281264 96784
rect 281316 96772 281322 96824
rect 282362 96772 282368 96824
rect 282420 96812 282426 96824
rect 282546 96812 282552 96824
rect 282420 96784 282552 96812
rect 282420 96772 282426 96784
rect 282546 96772 282552 96784
rect 282604 96772 282610 96824
rect 283558 96772 283564 96824
rect 283616 96812 283622 96824
rect 284018 96812 284024 96824
rect 283616 96784 284024 96812
rect 283616 96772 283622 96784
rect 284018 96772 284024 96784
rect 284076 96772 284082 96824
rect 286502 96772 286508 96824
rect 286560 96812 286566 96824
rect 286778 96812 286784 96824
rect 286560 96784 286784 96812
rect 286560 96772 286566 96784
rect 286778 96772 286784 96784
rect 286836 96772 286842 96824
rect 277578 96704 277584 96756
rect 277636 96744 277642 96756
rect 278590 96744 278596 96756
rect 277636 96716 278596 96744
rect 277636 96704 277642 96716
rect 278590 96704 278596 96716
rect 278648 96704 278654 96756
rect 279510 96704 279516 96756
rect 279568 96744 279574 96756
rect 287026 96744 287054 96852
rect 307018 96840 307024 96852
rect 307076 96840 307082 96892
rect 287146 96772 287152 96824
rect 287204 96812 287210 96824
rect 287790 96812 287796 96824
rect 287204 96784 287796 96812
rect 287204 96772 287210 96784
rect 287790 96772 287796 96784
rect 287848 96772 287854 96824
rect 289170 96772 289176 96824
rect 289228 96812 289234 96824
rect 289722 96812 289728 96824
rect 289228 96784 289728 96812
rect 289228 96772 289234 96784
rect 289722 96772 289728 96784
rect 289780 96772 289786 96824
rect 290734 96772 290740 96824
rect 290792 96812 290798 96824
rect 290918 96812 290924 96824
rect 290792 96784 290924 96812
rect 290792 96772 290798 96784
rect 290918 96772 290924 96784
rect 290976 96772 290982 96824
rect 291286 96772 291292 96824
rect 291344 96812 291350 96824
rect 291930 96812 291936 96824
rect 291344 96784 291936 96812
rect 291344 96772 291350 96784
rect 291930 96772 291936 96784
rect 291988 96772 291994 96824
rect 292206 96772 292212 96824
rect 292264 96812 292270 96824
rect 292482 96812 292488 96824
rect 292264 96784 292488 96812
rect 292264 96772 292270 96784
rect 292482 96772 292488 96784
rect 292540 96772 292546 96824
rect 294414 96772 294420 96824
rect 294472 96812 294478 96824
rect 295242 96812 295248 96824
rect 294472 96784 295248 96812
rect 294472 96772 294478 96784
rect 295242 96772 295248 96784
rect 295300 96772 295306 96824
rect 295518 96772 295524 96824
rect 295576 96812 295582 96824
rect 296438 96812 296444 96824
rect 295576 96784 296444 96812
rect 295576 96772 295582 96784
rect 296438 96772 296444 96784
rect 296496 96772 296502 96824
rect 296714 96772 296720 96824
rect 296772 96812 296778 96824
rect 298094 96812 298100 96824
rect 296772 96784 298100 96812
rect 296772 96772 296778 96784
rect 298094 96772 298100 96784
rect 298152 96772 298158 96824
rect 298186 96772 298192 96824
rect 298244 96812 298250 96824
rect 304350 96812 304356 96824
rect 298244 96784 304356 96812
rect 298244 96772 298250 96784
rect 304350 96772 304356 96784
rect 304408 96772 304414 96824
rect 279568 96716 287054 96744
rect 279568 96704 279574 96716
rect 287698 96704 287704 96756
rect 287756 96744 287762 96756
rect 288066 96744 288072 96756
rect 287756 96716 288072 96744
rect 287756 96704 287762 96716
rect 288066 96704 288072 96716
rect 288124 96704 288130 96756
rect 288526 96704 288532 96756
rect 288584 96744 288590 96756
rect 289538 96744 289544 96756
rect 288584 96716 289544 96744
rect 288584 96704 288590 96716
rect 289538 96704 289544 96716
rect 289596 96704 289602 96756
rect 291470 96704 291476 96756
rect 291528 96744 291534 96756
rect 292114 96744 292120 96756
rect 291528 96716 292120 96744
rect 291528 96704 291534 96716
rect 292114 96704 292120 96716
rect 292172 96704 292178 96756
rect 294506 96704 294512 96756
rect 294564 96744 294570 96756
rect 294966 96744 294972 96756
rect 294564 96716 294972 96744
rect 294564 96704 294570 96716
rect 294966 96704 294972 96716
rect 295024 96704 295030 96756
rect 296070 96704 296076 96756
rect 296128 96744 296134 96756
rect 296346 96744 296352 96756
rect 296128 96716 296352 96744
rect 296128 96704 296134 96716
rect 296346 96704 296352 96716
rect 296404 96704 296410 96756
rect 296990 96704 296996 96756
rect 297048 96744 297054 96756
rect 297818 96744 297824 96756
rect 297048 96716 297824 96744
rect 297048 96704 297054 96716
rect 297818 96704 297824 96716
rect 297876 96704 297882 96756
rect 298002 96704 298008 96756
rect 298060 96744 298066 96756
rect 304258 96744 304264 96756
rect 298060 96716 304264 96744
rect 298060 96704 298066 96716
rect 304258 96704 304264 96716
rect 304316 96704 304322 96756
rect 282730 96676 282736 96688
rect 277504 96648 282736 96676
rect 282730 96636 282736 96648
rect 282788 96636 282794 96688
rect 283098 96636 283104 96688
rect 283156 96676 283162 96688
rect 283834 96676 283840 96688
rect 283156 96648 283840 96676
rect 283156 96636 283162 96648
rect 283834 96636 283840 96648
rect 283892 96636 283898 96688
rect 287330 96636 287336 96688
rect 287388 96676 287394 96688
rect 287882 96676 287888 96688
rect 287388 96648 287888 96676
rect 287388 96636 287394 96648
rect 287882 96636 287888 96648
rect 287940 96636 287946 96688
rect 291838 96636 291844 96688
rect 291896 96676 291902 96688
rect 292298 96676 292304 96688
rect 291896 96648 292304 96676
rect 291896 96636 291902 96648
rect 292298 96636 292304 96648
rect 292356 96636 292362 96688
rect 294138 96636 294144 96688
rect 294196 96676 294202 96688
rect 294782 96676 294788 96688
rect 294196 96648 294788 96676
rect 294196 96636 294202 96648
rect 294782 96636 294788 96648
rect 294840 96636 294846 96688
rect 294874 96636 294880 96688
rect 294932 96676 294938 96688
rect 295150 96676 295156 96688
rect 294932 96648 295156 96676
rect 294932 96636 294938 96648
rect 295150 96636 295156 96648
rect 295208 96636 295214 96688
rect 295702 96636 295708 96688
rect 295760 96676 295766 96688
rect 296162 96676 296168 96688
rect 295760 96648 296168 96676
rect 295760 96636 295766 96648
rect 296162 96636 296168 96648
rect 296220 96636 296226 96688
rect 297266 96636 297272 96688
rect 297324 96676 297330 96688
rect 297910 96676 297916 96688
rect 297324 96648 297916 96676
rect 297324 96636 297330 96648
rect 297910 96636 297916 96648
rect 297968 96636 297974 96688
rect 324958 96608 324964 96620
rect 277366 96580 324964 96608
rect 274358 96500 274364 96552
rect 274416 96500 274422 96552
rect 275830 96500 275836 96552
rect 275888 96500 275894 96552
rect 277366 96472 277394 96580
rect 324958 96568 324964 96580
rect 325016 96568 325022 96620
rect 285582 96500 285588 96552
rect 285640 96540 285646 96552
rect 461578 96540 461584 96552
rect 285640 96512 461584 96540
rect 285640 96500 285646 96512
rect 461578 96500 461584 96512
rect 461636 96500 461642 96552
rect 258046 96444 277394 96472
rect 283742 96432 283748 96484
rect 283800 96472 283806 96484
rect 468478 96472 468484 96484
rect 283800 96444 468484 96472
rect 283800 96432 283806 96444
rect 468478 96432 468484 96444
rect 468536 96432 468542 96484
rect 179322 96364 179328 96416
rect 179380 96404 179386 96416
rect 230106 96404 230112 96416
rect 179380 96376 230112 96404
rect 179380 96364 179386 96376
rect 230106 96364 230112 96376
rect 230164 96364 230170 96416
rect 285030 96364 285036 96416
rect 285088 96404 285094 96416
rect 285398 96404 285404 96416
rect 285088 96376 285404 96404
rect 285088 96364 285094 96376
rect 285398 96364 285404 96376
rect 285456 96364 285462 96416
rect 472618 96404 472624 96416
rect 285508 96376 472624 96404
rect 176562 96296 176568 96348
rect 176620 96336 176626 96348
rect 227714 96336 227720 96348
rect 176620 96308 227720 96336
rect 176620 96296 176626 96308
rect 227714 96296 227720 96308
rect 227772 96296 227778 96348
rect 282822 96296 282828 96348
rect 282880 96336 282886 96348
rect 285508 96336 285536 96376
rect 472618 96364 472624 96376
rect 472676 96364 472682 96416
rect 475378 96336 475384 96348
rect 282880 96308 285536 96336
rect 285692 96308 475384 96336
rect 282880 96296 282886 96308
rect 173158 96228 173164 96280
rect 173216 96268 173222 96280
rect 228910 96268 228916 96280
rect 173216 96240 228916 96268
rect 173216 96228 173222 96240
rect 228910 96228 228916 96240
rect 228968 96228 228974 96280
rect 282086 96228 282092 96280
rect 282144 96268 282150 96280
rect 285692 96268 285720 96308
rect 475378 96296 475384 96308
rect 475436 96296 475442 96348
rect 282144 96240 285720 96268
rect 282144 96228 282150 96240
rect 285858 96228 285864 96280
rect 285916 96268 285922 96280
rect 479518 96268 479524 96280
rect 285916 96240 479524 96268
rect 285916 96228 285922 96240
rect 479518 96228 479524 96240
rect 479576 96228 479582 96280
rect 169662 96160 169668 96212
rect 169720 96200 169726 96212
rect 228358 96200 228364 96212
rect 169720 96172 228364 96200
rect 169720 96160 169726 96172
rect 228358 96160 228364 96172
rect 228416 96160 228422 96212
rect 281534 96160 281540 96212
rect 281592 96200 281598 96212
rect 483014 96200 483020 96212
rect 281592 96172 483020 96200
rect 281592 96160 281598 96172
rect 483014 96160 483020 96172
rect 483072 96160 483078 96212
rect 155218 96092 155224 96144
rect 155276 96132 155282 96144
rect 225966 96132 225972 96144
rect 155276 96104 225972 96132
rect 155276 96092 155282 96104
rect 225966 96092 225972 96104
rect 226024 96092 226030 96144
rect 283374 96092 283380 96144
rect 283432 96132 283438 96144
rect 494054 96132 494060 96144
rect 283432 96104 494060 96132
rect 283432 96092 283438 96104
rect 494054 96092 494060 96104
rect 494112 96092 494118 96144
rect 133782 96024 133788 96076
rect 133840 96064 133846 96076
rect 215294 96064 215300 96076
rect 133840 96036 215300 96064
rect 133840 96024 133846 96036
rect 215294 96024 215300 96036
rect 215352 96024 215358 96076
rect 284570 96024 284576 96076
rect 284628 96064 284634 96076
rect 500954 96064 500960 96076
rect 284628 96036 500960 96064
rect 284628 96024 284634 96036
rect 500954 96024 500960 96036
rect 501012 96024 501018 96076
rect 70302 95956 70308 96008
rect 70360 95996 70366 96008
rect 211614 95996 211620 96008
rect 70360 95968 211620 95996
rect 70360 95956 70366 95968
rect 211614 95956 211620 95968
rect 211672 95956 211678 96008
rect 280982 95956 280988 96008
rect 281040 95996 281046 96008
rect 281040 95968 285720 95996
rect 281040 95956 281046 95968
rect 17862 95888 17868 95940
rect 17920 95928 17926 95940
rect 202874 95928 202880 95940
rect 17920 95900 202880 95928
rect 17920 95888 17926 95900
rect 202874 95888 202880 95900
rect 202932 95888 202938 95940
rect 202966 95888 202972 95940
rect 203024 95928 203030 95940
rect 203702 95928 203708 95940
rect 203024 95900 203708 95928
rect 203024 95888 203030 95900
rect 203702 95888 203708 95900
rect 203760 95888 203766 95940
rect 247678 95888 247684 95940
rect 247736 95928 247742 95940
rect 282178 95928 282184 95940
rect 247736 95900 282184 95928
rect 247736 95888 247742 95900
rect 282178 95888 282184 95900
rect 282236 95888 282242 95940
rect 285692 95928 285720 95968
rect 285766 95956 285772 96008
rect 285824 95996 285830 96008
rect 507854 95996 507860 96008
rect 285824 95968 507860 95996
rect 285824 95956 285830 95968
rect 507854 95956 507860 95968
rect 507912 95956 507918 96008
rect 285858 95928 285864 95940
rect 285692 95900 285864 95928
rect 285858 95888 285864 95900
rect 285916 95888 285922 95940
rect 297358 95888 297364 95940
rect 297416 95928 297422 95940
rect 518894 95928 518900 95940
rect 297416 95900 518900 95928
rect 297416 95888 297422 95900
rect 518894 95888 518900 95900
rect 518952 95888 518958 95940
rect 165522 95820 165528 95872
rect 165580 95860 165586 95872
rect 208118 95860 208124 95872
rect 165580 95832 208124 95860
rect 165580 95820 165586 95832
rect 208118 95820 208124 95832
rect 208176 95820 208182 95872
rect 253014 95820 253020 95872
rect 253072 95860 253078 95872
rect 312538 95860 312544 95872
rect 253072 95832 312544 95860
rect 253072 95820 253078 95832
rect 312538 95820 312544 95832
rect 312596 95820 312602 95872
rect 191098 95752 191104 95804
rect 191156 95792 191162 95804
rect 231946 95792 231952 95804
rect 191156 95764 231952 95792
rect 191156 95752 191162 95764
rect 231946 95752 231952 95764
rect 232004 95752 232010 95804
rect 252462 95752 252468 95804
rect 252520 95792 252526 95804
rect 309134 95792 309140 95804
rect 252520 95764 309140 95792
rect 252520 95752 252526 95764
rect 309134 95752 309140 95764
rect 309192 95752 309198 95804
rect 197262 95684 197268 95736
rect 197320 95724 197326 95736
rect 233142 95724 233148 95736
rect 197320 95696 233148 95724
rect 197320 95684 197326 95696
rect 233142 95684 233148 95696
rect 233200 95684 233206 95736
rect 242894 95684 242900 95736
rect 242952 95724 242958 95736
rect 250438 95724 250444 95736
rect 242952 95696 250444 95724
rect 242952 95684 242958 95696
rect 250438 95684 250444 95696
rect 250496 95684 250502 95736
rect 251082 95684 251088 95736
rect 251140 95724 251146 95736
rect 302234 95724 302240 95736
rect 251140 95696 302240 95724
rect 251140 95684 251146 95696
rect 302234 95684 302240 95696
rect 302292 95684 302298 95736
rect 200022 95616 200028 95668
rect 200080 95656 200086 95668
rect 233878 95656 233884 95668
rect 200080 95628 233884 95656
rect 200080 95616 200086 95628
rect 233878 95616 233884 95628
rect 233936 95616 233942 95668
rect 256694 95616 256700 95668
rect 256752 95656 256758 95668
rect 306374 95656 306380 95668
rect 256752 95628 306380 95656
rect 256752 95616 256758 95628
rect 306374 95616 306380 95628
rect 306432 95616 306438 95668
rect 194502 95548 194508 95600
rect 194560 95588 194566 95600
rect 218054 95588 218060 95600
rect 194560 95560 218060 95588
rect 194560 95548 194566 95560
rect 218054 95548 218060 95560
rect 218112 95548 218118 95600
rect 249886 95548 249892 95600
rect 249944 95588 249950 95600
rect 298186 95588 298192 95600
rect 249944 95560 298192 95588
rect 249944 95548 249950 95560
rect 298186 95548 298192 95560
rect 298244 95548 298250 95600
rect 262858 95480 262864 95532
rect 262916 95520 262922 95532
rect 299474 95520 299480 95532
rect 262916 95492 299480 95520
rect 262916 95480 262922 95492
rect 299474 95480 299480 95492
rect 299532 95480 299538 95532
rect 287514 95412 287520 95464
rect 287572 95452 287578 95464
rect 297358 95452 297364 95464
rect 287572 95424 297364 95452
rect 287572 95412 287578 95424
rect 297358 95412 297364 95424
rect 297416 95412 297422 95464
rect 233142 95344 233148 95396
rect 233200 95384 233206 95396
rect 239122 95384 239128 95396
rect 233200 95356 239128 95384
rect 233200 95344 233206 95356
rect 239122 95344 239128 95356
rect 239180 95344 239186 95396
rect 234430 95276 234436 95328
rect 234488 95316 234494 95328
rect 239950 95316 239956 95328
rect 234488 95288 239956 95316
rect 234488 95276 234494 95288
rect 239950 95276 239956 95288
rect 240008 95276 240014 95328
rect 228634 95208 228640 95260
rect 228692 95248 228698 95260
rect 233970 95248 233976 95260
rect 228692 95220 233976 95248
rect 228692 95208 228698 95220
rect 233970 95208 233976 95220
rect 234028 95208 234034 95260
rect 162762 95140 162768 95192
rect 162820 95180 162826 95192
rect 227346 95180 227352 95192
rect 162820 95152 227352 95180
rect 162820 95140 162826 95152
rect 227346 95140 227352 95152
rect 227404 95140 227410 95192
rect 286962 95140 286968 95192
rect 287020 95180 287026 95192
rect 454678 95180 454684 95192
rect 287020 95152 454684 95180
rect 287020 95140 287026 95152
rect 454678 95140 454684 95152
rect 454736 95140 454742 95192
rect 158622 95072 158628 95124
rect 158680 95112 158686 95124
rect 226518 95112 226524 95124
rect 158680 95084 226524 95112
rect 158680 95072 158686 95084
rect 226518 95072 226524 95084
rect 226576 95072 226582 95124
rect 279694 95072 279700 95124
rect 279752 95112 279758 95124
rect 464338 95112 464344 95124
rect 279752 95084 464344 95112
rect 279752 95072 279758 95084
rect 464338 95072 464344 95084
rect 464396 95072 464402 95124
rect 144822 95004 144828 95056
rect 144880 95044 144886 95056
rect 212534 95044 212540 95056
rect 144880 95016 212540 95044
rect 144880 95004 144886 95016
rect 212534 95004 212540 95016
rect 212592 95004 212598 95056
rect 292390 95004 292396 95056
rect 292448 95044 292454 95056
rect 485038 95044 485044 95056
rect 292448 95016 485044 95044
rect 292448 95004 292454 95016
rect 485038 95004 485044 95016
rect 485096 95004 485102 95056
rect 147582 94936 147588 94988
rect 147640 94976 147646 94988
rect 224770 94976 224776 94988
rect 147640 94948 224776 94976
rect 147640 94936 147646 94948
rect 224770 94936 224776 94948
rect 224828 94936 224834 94988
rect 291102 94936 291108 94988
rect 291160 94976 291166 94988
rect 489178 94976 489184 94988
rect 291160 94948 489184 94976
rect 291160 94936 291166 94948
rect 489178 94936 489184 94948
rect 489236 94936 489242 94988
rect 137278 94868 137284 94920
rect 137336 94908 137342 94920
rect 223022 94908 223028 94920
rect 137336 94880 223028 94908
rect 137336 94868 137342 94880
rect 223022 94868 223028 94880
rect 223080 94868 223086 94920
rect 289630 94868 289636 94920
rect 289688 94908 289694 94920
rect 502978 94908 502984 94920
rect 289688 94880 502984 94908
rect 289688 94868 289694 94880
rect 502978 94868 502984 94880
rect 503036 94868 503042 94920
rect 128262 94800 128268 94852
rect 128320 94840 128326 94852
rect 221366 94840 221372 94852
rect 128320 94812 221372 94840
rect 128320 94800 128326 94812
rect 221366 94800 221372 94812
rect 221424 94800 221430 94852
rect 286318 94800 286324 94852
rect 286376 94840 286382 94852
rect 511994 94840 512000 94852
rect 286376 94812 512000 94840
rect 286376 94800 286382 94812
rect 511994 94800 512000 94812
rect 512052 94800 512058 94852
rect 78582 94732 78588 94784
rect 78640 94772 78646 94784
rect 213086 94772 213092 94784
rect 78640 94744 213092 94772
rect 78640 94732 78646 94744
rect 213086 94732 213092 94744
rect 213144 94732 213150 94784
rect 288158 94732 288164 94784
rect 288216 94772 288222 94784
rect 520918 94772 520924 94784
rect 288216 94744 520924 94772
rect 288216 94732 288222 94744
rect 520918 94732 520924 94744
rect 520976 94732 520982 94784
rect 64782 94664 64788 94716
rect 64840 94704 64846 94716
rect 210786 94704 210792 94716
rect 64840 94676 210792 94704
rect 64840 94664 64846 94676
rect 210786 94664 210792 94676
rect 210844 94664 210850 94716
rect 229738 94664 229744 94716
rect 229796 94704 229802 94716
rect 237558 94704 237564 94716
rect 229796 94676 237564 94704
rect 229796 94664 229802 94676
rect 237558 94664 237564 94676
rect 237616 94664 237622 94716
rect 288710 94664 288716 94716
rect 288768 94704 288774 94716
rect 525794 94704 525800 94716
rect 288768 94676 525800 94704
rect 288768 94664 288774 94676
rect 525794 94664 525800 94676
rect 525852 94664 525858 94716
rect 37090 94596 37096 94648
rect 37148 94636 37154 94648
rect 206278 94636 206284 94648
rect 37148 94608 206284 94636
rect 37148 94596 37154 94608
rect 206278 94596 206284 94608
rect 206336 94596 206342 94648
rect 244918 94596 244924 94648
rect 244976 94636 244982 94648
rect 262858 94636 262864 94648
rect 244976 94608 262864 94636
rect 244976 94596 244982 94608
rect 262858 94596 262864 94608
rect 262916 94596 262922 94648
rect 290550 94596 290556 94648
rect 290608 94636 290614 94648
rect 536834 94636 536840 94648
rect 290608 94608 536840 94636
rect 290608 94596 290614 94608
rect 536834 94596 536840 94608
rect 536892 94596 536898 94648
rect 33778 94528 33784 94580
rect 33836 94568 33842 94580
rect 205266 94568 205272 94580
rect 33836 94540 205272 94568
rect 33836 94528 33842 94540
rect 205266 94528 205272 94540
rect 205324 94528 205330 94580
rect 208578 94528 208584 94580
rect 208636 94568 208642 94580
rect 209498 94568 209504 94580
rect 208636 94540 209504 94568
rect 208636 94528 208642 94540
rect 209498 94528 209504 94540
rect 209556 94528 209562 94580
rect 210142 94528 210148 94580
rect 210200 94568 210206 94580
rect 210602 94568 210608 94580
rect 210200 94540 210608 94568
rect 210200 94528 210206 94540
rect 210602 94528 210608 94540
rect 210660 94528 210666 94580
rect 212902 94528 212908 94580
rect 212960 94568 212966 94580
rect 213546 94568 213552 94580
rect 212960 94540 213552 94568
rect 212960 94528 212966 94540
rect 213546 94528 213552 94540
rect 213604 94528 213610 94580
rect 214098 94528 214104 94580
rect 214156 94568 214162 94580
rect 214742 94568 214748 94580
rect 214156 94540 214748 94568
rect 214156 94528 214162 94540
rect 214742 94528 214748 94540
rect 214800 94528 214806 94580
rect 233602 94528 233608 94580
rect 233660 94568 233666 94580
rect 234246 94568 234252 94580
rect 233660 94540 234252 94568
rect 233660 94528 233666 94540
rect 234246 94528 234252 94540
rect 234304 94528 234310 94580
rect 248046 94528 248052 94580
rect 248104 94568 248110 94580
rect 285674 94568 285680 94580
rect 248104 94540 285680 94568
rect 248104 94528 248110 94540
rect 285674 94528 285680 94540
rect 285732 94528 285738 94580
rect 291746 94528 291752 94580
rect 291804 94568 291810 94580
rect 543734 94568 543740 94580
rect 291804 94540 543740 94568
rect 291804 94528 291810 94540
rect 543734 94528 543740 94540
rect 543792 94528 543798 94580
rect 25498 94460 25504 94512
rect 25556 94500 25562 94512
rect 203610 94500 203616 94512
rect 25556 94472 203616 94500
rect 25556 94460 25562 94472
rect 203610 94460 203616 94472
rect 203668 94460 203674 94512
rect 209958 94460 209964 94512
rect 210016 94500 210022 94512
rect 210878 94500 210884 94512
rect 210016 94472 210884 94500
rect 210016 94460 210022 94472
rect 210878 94460 210884 94472
rect 210936 94460 210942 94512
rect 224862 94460 224868 94512
rect 224920 94500 224926 94512
rect 231854 94500 231860 94512
rect 224920 94472 231860 94500
rect 224920 94460 224926 94472
rect 231854 94460 231860 94472
rect 231912 94460 231918 94512
rect 249702 94460 249708 94512
rect 249760 94500 249766 94512
rect 293218 94500 293224 94512
rect 249760 94472 293224 94500
rect 249760 94460 249766 94472
rect 293218 94460 293224 94472
rect 293276 94460 293282 94512
rect 293402 94460 293408 94512
rect 293460 94500 293466 94512
rect 293770 94500 293776 94512
rect 293460 94472 293776 94500
rect 293460 94460 293466 94472
rect 293770 94460 293776 94472
rect 293828 94460 293834 94512
rect 295334 94460 295340 94512
rect 295392 94500 295398 94512
rect 558178 94500 558184 94512
rect 295392 94472 558184 94500
rect 295392 94460 295398 94472
rect 558178 94460 558184 94472
rect 558236 94460 558242 94512
rect 166902 94392 166908 94444
rect 166960 94432 166966 94444
rect 227990 94432 227996 94444
rect 166960 94404 227996 94432
rect 166960 94392 166966 94404
rect 227990 94392 227996 94404
rect 228048 94392 228054 94444
rect 230842 94392 230848 94444
rect 230900 94432 230906 94444
rect 231670 94432 231676 94444
rect 230900 94404 231676 94432
rect 230900 94392 230906 94404
rect 231670 94392 231676 94404
rect 231728 94392 231734 94444
rect 259822 94392 259828 94444
rect 259880 94432 259886 94444
rect 353938 94432 353944 94444
rect 259880 94404 353944 94432
rect 259880 94392 259886 94404
rect 353938 94392 353944 94404
rect 353996 94392 354002 94444
rect 157242 94324 157248 94376
rect 157300 94364 157306 94376
rect 216674 94364 216680 94376
rect 157300 94336 216680 94364
rect 157300 94324 157306 94336
rect 216674 94324 216680 94336
rect 216732 94324 216738 94376
rect 231118 94324 231124 94376
rect 231176 94364 231182 94376
rect 236914 94364 236920 94376
rect 231176 94336 236920 94364
rect 231176 94324 231182 94336
rect 236914 94324 236920 94336
rect 236972 94324 236978 94376
rect 255866 94324 255872 94376
rect 255924 94364 255930 94376
rect 331214 94364 331220 94376
rect 255924 94336 331220 94364
rect 255924 94324 255930 94336
rect 331214 94324 331220 94336
rect 331272 94324 331278 94376
rect 174538 94256 174544 94308
rect 174596 94296 174602 94308
rect 229186 94296 229192 94308
rect 174596 94268 229192 94296
rect 174596 94256 174602 94268
rect 229186 94256 229192 94268
rect 229244 94256 229250 94308
rect 253750 94256 253756 94308
rect 253808 94296 253814 94308
rect 316034 94296 316040 94308
rect 253808 94268 316040 94296
rect 253808 94256 253814 94268
rect 316034 94256 316040 94268
rect 316092 94256 316098 94308
rect 177942 94188 177948 94240
rect 178000 94228 178006 94240
rect 229646 94228 229652 94240
rect 178000 94200 229652 94228
rect 178000 94188 178006 94200
rect 229646 94188 229652 94200
rect 229704 94188 229710 94240
rect 252830 94188 252836 94240
rect 252888 94228 252894 94240
rect 313274 94228 313280 94240
rect 252888 94200 313280 94228
rect 252888 94188 252894 94200
rect 313274 94188 313280 94200
rect 313332 94188 313338 94240
rect 184842 94120 184848 94172
rect 184900 94160 184906 94172
rect 230750 94160 230756 94172
rect 184900 94132 230756 94160
rect 184900 94120 184906 94132
rect 230750 94120 230756 94132
rect 230808 94120 230814 94172
rect 262766 94120 262772 94172
rect 262824 94160 262830 94172
rect 320174 94160 320180 94172
rect 262824 94132 320180 94160
rect 262824 94120 262830 94132
rect 320174 94120 320180 94132
rect 320232 94120 320238 94172
rect 198642 94052 198648 94104
rect 198700 94092 198706 94104
rect 233234 94092 233240 94104
rect 198700 94064 233240 94092
rect 198700 94052 198706 94064
rect 233234 94052 233240 94064
rect 233292 94052 233298 94104
rect 292666 94052 292672 94104
rect 292724 94092 292730 94104
rect 293678 94092 293684 94104
rect 292724 94064 293684 94092
rect 292724 94052 292730 94064
rect 293678 94052 293684 94064
rect 293736 94052 293742 94104
rect 160002 93780 160008 93832
rect 160060 93820 160066 93832
rect 226794 93820 226800 93832
rect 160060 93792 226800 93820
rect 160060 93780 160066 93792
rect 226794 93780 226800 93792
rect 226852 93780 226858 93832
rect 261846 93780 261852 93832
rect 261904 93820 261910 93832
rect 360838 93820 360844 93832
rect 261904 93792 360844 93820
rect 261904 93780 261910 93792
rect 360838 93780 360844 93792
rect 360896 93780 360902 93832
rect 155862 93712 155868 93764
rect 155920 93752 155926 93764
rect 226058 93752 226064 93764
rect 155920 93724 226064 93752
rect 155920 93712 155926 93724
rect 226058 93712 226064 93724
rect 226116 93712 226122 93764
rect 262122 93712 262128 93764
rect 262180 93752 262186 93764
rect 364978 93752 364984 93764
rect 262180 93724 364984 93752
rect 262180 93712 262186 93724
rect 364978 93712 364984 93724
rect 365036 93712 365042 93764
rect 148962 93644 148968 93696
rect 149020 93684 149026 93696
rect 218790 93684 218796 93696
rect 149020 93656 218796 93684
rect 149020 93644 149026 93656
rect 218790 93644 218796 93656
rect 218848 93644 218854 93696
rect 263318 93644 263324 93696
rect 263376 93684 263382 93696
rect 367738 93684 367744 93696
rect 263376 93656 367744 93684
rect 263376 93644 263382 93656
rect 367738 93644 367744 93656
rect 367796 93644 367802 93696
rect 153102 93576 153108 93628
rect 153160 93616 153166 93628
rect 225414 93616 225420 93628
rect 153160 93588 225420 93616
rect 153160 93576 153166 93588
rect 225414 93576 225420 93588
rect 225472 93576 225478 93628
rect 264790 93576 264796 93628
rect 264848 93616 264854 93628
rect 374638 93616 374644 93628
rect 264848 93588 374644 93616
rect 264848 93576 264854 93588
rect 374638 93576 374644 93588
rect 374696 93576 374702 93628
rect 144730 93508 144736 93560
rect 144788 93548 144794 93560
rect 224034 93548 224040 93560
rect 144788 93520 224040 93548
rect 144788 93508 144794 93520
rect 224034 93508 224040 93520
rect 224092 93508 224098 93560
rect 270402 93508 270408 93560
rect 270460 93548 270466 93560
rect 416774 93548 416780 93560
rect 270460 93520 416780 93548
rect 270460 93508 270466 93520
rect 416774 93508 416780 93520
rect 416832 93508 416838 93560
rect 142062 93440 142068 93492
rect 142120 93480 142126 93492
rect 223666 93480 223672 93492
rect 142120 93452 223672 93480
rect 142120 93440 142126 93452
rect 223666 93440 223672 93452
rect 223724 93440 223730 93492
rect 273162 93440 273168 93492
rect 273220 93480 273226 93492
rect 421558 93480 421564 93492
rect 273220 93452 421564 93480
rect 273220 93440 273226 93452
rect 421558 93440 421564 93452
rect 421616 93440 421622 93492
rect 131022 93372 131028 93424
rect 131080 93412 131086 93424
rect 221458 93412 221464 93424
rect 131080 93384 221464 93412
rect 131080 93372 131086 93384
rect 221458 93372 221464 93384
rect 221516 93372 221522 93424
rect 275922 93372 275928 93424
rect 275980 93412 275986 93424
rect 448514 93412 448520 93424
rect 275980 93384 448520 93412
rect 275980 93372 275986 93384
rect 448514 93372 448520 93384
rect 448572 93372 448578 93424
rect 84102 93304 84108 93356
rect 84160 93344 84166 93356
rect 213822 93344 213828 93356
rect 84160 93316 213828 93344
rect 84160 93304 84166 93316
rect 213822 93304 213828 93316
rect 213880 93304 213886 93356
rect 293494 93304 293500 93356
rect 293552 93344 293558 93356
rect 554038 93344 554044 93356
rect 293552 93316 554044 93344
rect 293552 93304 293558 93316
rect 554038 93304 554044 93316
rect 554096 93304 554102 93356
rect 73062 93236 73068 93288
rect 73120 93276 73126 93288
rect 212074 93276 212080 93288
rect 73120 93248 212080 93276
rect 73120 93236 73126 93248
rect 212074 93236 212080 93248
rect 212132 93236 212138 93288
rect 294690 93236 294696 93288
rect 294748 93276 294754 93288
rect 561674 93276 561680 93288
rect 294748 93248 561680 93276
rect 294748 93236 294754 93248
rect 561674 93236 561680 93248
rect 561732 93236 561738 93288
rect 68278 93168 68284 93220
rect 68336 93208 68342 93220
rect 210050 93208 210056 93220
rect 68336 93180 210056 93208
rect 68336 93168 68342 93180
rect 210050 93168 210056 93180
rect 210108 93168 210114 93220
rect 243630 93168 243636 93220
rect 243688 93208 243694 93220
rect 257338 93208 257344 93220
rect 243688 93180 257344 93208
rect 243688 93168 243694 93180
rect 257338 93168 257344 93180
rect 257396 93168 257402 93220
rect 295978 93168 295984 93220
rect 296036 93208 296042 93220
rect 568574 93208 568580 93220
rect 296036 93180 568580 93208
rect 296036 93168 296042 93180
rect 568574 93168 568580 93180
rect 568632 93168 568638 93220
rect 14458 93100 14464 93152
rect 14516 93140 14522 93152
rect 201494 93140 201500 93152
rect 14516 93112 201500 93140
rect 14516 93100 14522 93112
rect 201494 93100 201500 93112
rect 201552 93100 201558 93152
rect 246850 93100 246856 93152
rect 246908 93140 246914 93152
rect 261478 93140 261484 93152
rect 246908 93112 261484 93140
rect 246908 93100 246914 93112
rect 261478 93100 261484 93112
rect 261536 93100 261542 93152
rect 296530 93100 296536 93152
rect 296588 93140 296594 93152
rect 572714 93140 572720 93152
rect 296588 93112 572720 93140
rect 296588 93100 296594 93112
rect 572714 93100 572720 93112
rect 572772 93100 572778 93152
rect 170398 93032 170404 93084
rect 170456 93072 170462 93084
rect 228450 93072 228456 93084
rect 170456 93044 228456 93072
rect 170456 93032 170462 93044
rect 228450 93032 228456 93044
rect 228508 93032 228514 93084
rect 257982 93032 257988 93084
rect 258040 93072 258046 93084
rect 340874 93072 340880 93084
rect 258040 93044 340880 93072
rect 258040 93032 258046 93044
rect 340874 93032 340880 93044
rect 340932 93032 340938 93084
rect 180702 92964 180708 93016
rect 180760 93004 180766 93016
rect 230198 93004 230204 93016
rect 180760 92976 230204 93004
rect 180760 92964 180766 92976
rect 230198 92964 230204 92976
rect 230256 92964 230262 93016
rect 257798 92964 257804 93016
rect 257856 93004 257862 93016
rect 338114 93004 338120 93016
rect 257856 92976 338120 93004
rect 257856 92964 257862 92976
rect 338114 92964 338120 92976
rect 338172 92964 338178 93016
rect 188338 92896 188344 92948
rect 188396 92936 188402 92948
rect 231394 92936 231400 92948
rect 188396 92908 231400 92936
rect 188396 92896 188402 92908
rect 231394 92896 231400 92908
rect 231452 92896 231458 92948
rect 256510 92896 256516 92948
rect 256568 92936 256574 92948
rect 333974 92936 333980 92948
rect 256568 92908 333980 92936
rect 256568 92896 256574 92908
rect 333974 92896 333980 92908
rect 334032 92896 334038 92948
rect 229830 92556 229836 92608
rect 229888 92596 229894 92608
rect 236546 92596 236552 92608
rect 229888 92568 236552 92596
rect 229888 92556 229894 92568
rect 236546 92556 236552 92568
rect 236604 92556 236610 92608
rect 231210 92488 231216 92540
rect 231268 92528 231274 92540
rect 234614 92528 234620 92540
rect 231268 92500 234620 92528
rect 231268 92488 231274 92500
rect 234614 92488 234620 92500
rect 234672 92488 234678 92540
rect 177850 92420 177856 92472
rect 177908 92460 177914 92472
rect 229922 92460 229928 92472
rect 177908 92432 229928 92460
rect 177908 92420 177914 92432
rect 229922 92420 229928 92432
rect 229980 92420 229986 92472
rect 264882 92420 264888 92472
rect 264940 92460 264946 92472
rect 378778 92460 378784 92472
rect 264940 92432 378784 92460
rect 264940 92420 264946 92432
rect 378778 92420 378784 92432
rect 378836 92420 378842 92472
rect 175182 92352 175188 92404
rect 175240 92392 175246 92404
rect 229370 92392 229376 92404
rect 175240 92364 229376 92392
rect 175240 92352 175246 92364
rect 229370 92352 229376 92364
rect 229428 92352 229434 92404
rect 264606 92352 264612 92404
rect 264664 92392 264670 92404
rect 382918 92392 382924 92404
rect 264664 92364 382924 92392
rect 264664 92352 264670 92364
rect 382918 92352 382924 92364
rect 382976 92352 382982 92404
rect 169018 92284 169024 92336
rect 169076 92324 169082 92336
rect 228174 92324 228180 92336
rect 169076 92296 228180 92324
rect 169076 92284 169082 92296
rect 228174 92284 228180 92296
rect 228232 92284 228238 92336
rect 266998 92284 267004 92336
rect 267056 92324 267062 92336
rect 387794 92324 387800 92336
rect 267056 92296 387800 92324
rect 267056 92284 267062 92296
rect 387794 92284 387800 92296
rect 387852 92284 387858 92336
rect 164142 92216 164148 92268
rect 164200 92256 164206 92268
rect 227438 92256 227444 92268
rect 164200 92228 227444 92256
rect 164200 92216 164206 92228
rect 227438 92216 227444 92228
rect 227496 92216 227502 92268
rect 266262 92216 266268 92268
rect 266320 92256 266326 92268
rect 389818 92256 389824 92268
rect 266320 92228 389824 92256
rect 266320 92216 266326 92228
rect 389818 92216 389824 92228
rect 389876 92216 389882 92268
rect 128170 92148 128176 92200
rect 128228 92188 128234 92200
rect 221550 92188 221556 92200
rect 128228 92160 221556 92188
rect 128228 92148 128234 92160
rect 221550 92148 221556 92160
rect 221608 92148 221614 92200
rect 272886 92148 272892 92200
rect 272944 92188 272950 92200
rect 430574 92188 430580 92200
rect 272944 92160 430580 92188
rect 272944 92148 272950 92160
rect 430574 92148 430580 92160
rect 430632 92148 430638 92200
rect 104158 92080 104164 92132
rect 104216 92120 104222 92132
rect 217042 92120 217048 92132
rect 104216 92092 217048 92120
rect 104216 92080 104222 92092
rect 217042 92080 217048 92092
rect 217100 92080 217106 92132
rect 272978 92080 272984 92132
rect 273036 92120 273042 92132
rect 432598 92120 432604 92132
rect 273036 92092 432604 92120
rect 273036 92080 273042 92092
rect 432598 92080 432604 92092
rect 432656 92080 432662 92132
rect 79962 92012 79968 92064
rect 80020 92052 80026 92064
rect 213270 92052 213276 92064
rect 80020 92024 213276 92052
rect 80020 92012 80026 92024
rect 213270 92012 213276 92024
rect 213328 92012 213334 92064
rect 277302 92012 277308 92064
rect 277360 92052 277366 92064
rect 446398 92052 446404 92064
rect 277360 92024 446404 92052
rect 277360 92012 277366 92024
rect 446398 92012 446404 92024
rect 446456 92012 446462 92064
rect 77202 91944 77208 91996
rect 77260 91984 77266 91996
rect 212810 91984 212816 91996
rect 77260 91956 212816 91984
rect 77260 91944 77266 91956
rect 212810 91944 212816 91956
rect 212868 91944 212874 91996
rect 277026 91944 277032 91996
rect 277084 91984 277090 91996
rect 453298 91984 453304 91996
rect 277084 91956 453304 91984
rect 277084 91944 277090 91956
rect 453298 91944 453304 91956
rect 453356 91944 453362 91996
rect 54478 91876 54484 91928
rect 54536 91916 54542 91928
rect 208486 91916 208492 91928
rect 54536 91888 208492 91916
rect 54536 91876 54542 91888
rect 208486 91876 208492 91888
rect 208544 91876 208550 91928
rect 278682 91876 278688 91928
rect 278740 91916 278746 91928
rect 460198 91916 460204 91928
rect 278740 91888 460204 91916
rect 278740 91876 278746 91888
rect 460198 91876 460204 91888
rect 460256 91876 460262 91928
rect 45462 91808 45468 91860
rect 45520 91848 45526 91860
rect 207474 91848 207480 91860
rect 45520 91820 207480 91848
rect 45520 91808 45526 91820
rect 207474 91808 207480 91820
rect 207532 91808 207538 91860
rect 246942 91808 246948 91860
rect 247000 91848 247006 91860
rect 264238 91848 264244 91860
rect 247000 91820 264244 91848
rect 247000 91808 247006 91820
rect 264238 91808 264244 91820
rect 264296 91808 264302 91860
rect 279878 91808 279884 91860
rect 279936 91848 279942 91860
rect 465718 91848 465724 91860
rect 279936 91820 465724 91848
rect 279936 91808 279942 91820
rect 465718 91808 465724 91820
rect 465776 91808 465782 91860
rect 23382 91740 23388 91792
rect 23440 91780 23446 91792
rect 202966 91780 202972 91792
rect 23440 91752 202972 91780
rect 23440 91740 23446 91752
rect 202966 91740 202972 91752
rect 203024 91740 203030 91792
rect 230382 91740 230388 91792
rect 230440 91780 230446 91792
rect 239398 91780 239404 91792
rect 230440 91752 239404 91780
rect 230440 91740 230446 91752
rect 239398 91740 239404 91752
rect 239456 91740 239462 91792
rect 243998 91740 244004 91792
rect 244056 91780 244062 91792
rect 262214 91780 262220 91792
rect 244056 91752 262220 91780
rect 244056 91740 244062 91752
rect 262214 91740 262220 91752
rect 262272 91740 262278 91792
rect 287790 91740 287796 91792
rect 287848 91780 287854 91792
rect 515398 91780 515404 91792
rect 287848 91752 515404 91780
rect 287848 91740 287854 91752
rect 515398 91740 515404 91752
rect 515456 91740 515462 91792
rect 182082 91672 182088 91724
rect 182140 91712 182146 91724
rect 230658 91712 230664 91724
rect 182140 91684 230664 91712
rect 182140 91672 182146 91684
rect 230658 91672 230664 91684
rect 230716 91672 230722 91724
rect 233418 91672 233424 91724
rect 233476 91712 233482 91724
rect 234062 91712 234068 91724
rect 233476 91684 234068 91712
rect 233476 91672 233482 91684
rect 234062 91672 234068 91684
rect 234120 91672 234126 91724
rect 260742 91672 260748 91724
rect 260800 91712 260806 91724
rect 353294 91712 353300 91724
rect 260800 91684 353300 91712
rect 260800 91672 260806 91684
rect 353294 91672 353300 91684
rect 353352 91672 353358 91724
rect 187050 91604 187056 91656
rect 187108 91644 187114 91656
rect 231026 91644 231032 91656
rect 187108 91616 231032 91644
rect 187108 91604 187114 91616
rect 231026 91604 231032 91616
rect 231084 91604 231090 91656
rect 256050 91604 256056 91656
rect 256108 91644 256114 91656
rect 328454 91644 328460 91656
rect 256108 91616 328460 91644
rect 256108 91604 256114 91616
rect 328454 91604 328460 91616
rect 328512 91604 328518 91656
rect 232222 90992 232228 91044
rect 232280 91032 232286 91044
rect 232590 91032 232596 91044
rect 232280 91004 232596 91032
rect 232280 90992 232286 91004
rect 232590 90992 232596 91004
rect 232648 90992 232654 91044
rect 274542 90992 274548 91044
rect 274600 91032 274606 91044
rect 407758 91032 407764 91044
rect 274600 91004 407764 91032
rect 274600 90992 274606 91004
rect 407758 90992 407764 91004
rect 407816 90992 407822 91044
rect 153010 90924 153016 90976
rect 153068 90964 153074 90976
rect 225690 90964 225696 90976
rect 153068 90936 225696 90964
rect 153068 90924 153074 90936
rect 225690 90924 225696 90936
rect 225748 90924 225754 90976
rect 269022 90924 269028 90976
rect 269080 90964 269086 90976
rect 403618 90964 403624 90976
rect 269080 90936 403624 90964
rect 269080 90924 269086 90936
rect 403618 90924 403624 90936
rect 403676 90924 403682 90976
rect 146202 90856 146208 90908
rect 146260 90896 146266 90908
rect 224494 90896 224500 90908
rect 146260 90868 224500 90896
rect 146260 90856 146266 90868
rect 224494 90856 224500 90868
rect 224552 90856 224558 90908
rect 289262 90856 289268 90908
rect 289320 90896 289326 90908
rect 471238 90896 471244 90908
rect 289320 90868 471244 90896
rect 289320 90856 289326 90868
rect 471238 90856 471244 90868
rect 471296 90856 471302 90908
rect 112438 90788 112444 90840
rect 112496 90828 112502 90840
rect 219066 90828 219072 90840
rect 112496 90800 219072 90828
rect 112496 90788 112502 90800
rect 219066 90788 219072 90800
rect 219124 90788 219130 90840
rect 278406 90788 278412 90840
rect 278464 90828 278470 90840
rect 465166 90828 465172 90840
rect 278464 90800 465172 90828
rect 278464 90788 278470 90800
rect 465166 90788 465172 90800
rect 465224 90788 465230 90840
rect 108942 90720 108948 90772
rect 109000 90760 109006 90772
rect 218882 90760 218888 90772
rect 109000 90732 218888 90760
rect 109000 90720 109006 90732
rect 218882 90720 218888 90732
rect 218940 90720 218946 90772
rect 282638 90720 282644 90772
rect 282696 90760 282702 90772
rect 476758 90760 476764 90772
rect 282696 90732 476764 90760
rect 282696 90720 282702 90732
rect 476758 90720 476764 90732
rect 476816 90720 476822 90772
rect 105538 90652 105544 90704
rect 105596 90692 105602 90704
rect 217502 90692 217508 90704
rect 105596 90664 217508 90692
rect 105596 90652 105602 90664
rect 217502 90652 217508 90664
rect 217560 90652 217566 90704
rect 282546 90652 282552 90704
rect 282604 90692 282610 90704
rect 486418 90692 486424 90704
rect 282604 90664 486424 90692
rect 282604 90652 282610 90664
rect 486418 90652 486424 90664
rect 486476 90652 486482 90704
rect 90358 90584 90364 90636
rect 90416 90624 90422 90636
rect 214926 90624 214932 90636
rect 90416 90596 214932 90624
rect 90416 90584 90422 90596
rect 214926 90584 214932 90596
rect 214984 90584 214990 90636
rect 284018 90584 284024 90636
rect 284076 90624 284082 90636
rect 493318 90624 493324 90636
rect 284076 90596 493324 90624
rect 284076 90584 284082 90596
rect 493318 90584 493324 90596
rect 493376 90584 493382 90636
rect 75178 90516 75184 90568
rect 75236 90556 75242 90568
rect 211338 90556 211344 90568
rect 75236 90528 211344 90556
rect 75236 90516 75242 90528
rect 211338 90516 211344 90528
rect 211396 90516 211402 90568
rect 283926 90516 283932 90568
rect 283984 90556 283990 90568
rect 497458 90556 497464 90568
rect 283984 90528 497464 90556
rect 283984 90516 283990 90528
rect 497458 90516 497464 90528
rect 497516 90516 497522 90568
rect 65518 90448 65524 90500
rect 65576 90488 65582 90500
rect 209314 90488 209320 90500
rect 65576 90460 209320 90488
rect 65576 90448 65582 90460
rect 209314 90448 209320 90460
rect 209372 90448 209378 90500
rect 285122 90448 285128 90500
rect 285180 90488 285186 90500
rect 500218 90488 500224 90500
rect 285180 90460 500224 90488
rect 285180 90448 285186 90460
rect 500218 90448 500224 90460
rect 500276 90448 500282 90500
rect 53098 90380 53104 90432
rect 53156 90420 53162 90432
rect 208026 90420 208032 90432
rect 53156 90392 208032 90420
rect 53156 90380 53162 90392
rect 208026 90380 208032 90392
rect 208084 90380 208090 90432
rect 286686 90380 286692 90432
rect 286744 90420 286750 90432
rect 504358 90420 504364 90432
rect 286744 90392 504364 90420
rect 286744 90380 286750 90392
rect 504358 90380 504364 90392
rect 504416 90380 504422 90432
rect 41322 90312 41328 90364
rect 41380 90352 41386 90364
rect 206738 90352 206744 90364
rect 41380 90324 206744 90352
rect 41380 90312 41386 90324
rect 206738 90312 206744 90324
rect 206796 90312 206802 90364
rect 217318 90312 217324 90364
rect 217376 90352 217382 90364
rect 234338 90352 234344 90364
rect 217376 90324 234344 90352
rect 217376 90312 217382 90324
rect 234338 90312 234344 90324
rect 234396 90312 234402 90364
rect 244090 90312 244096 90364
rect 244148 90352 244154 90364
rect 255958 90352 255964 90364
rect 244148 90324 255964 90352
rect 244148 90312 244154 90324
rect 255958 90312 255964 90324
rect 256016 90312 256022 90364
rect 291930 90312 291936 90364
rect 291988 90352 291994 90364
rect 540238 90352 540244 90364
rect 291988 90324 540244 90352
rect 291988 90312 291994 90324
rect 540238 90312 540244 90324
rect 540296 90312 540302 90364
rect 263410 90244 263416 90296
rect 263468 90284 263474 90296
rect 356698 90284 356704 90296
rect 263468 90256 356704 90284
rect 263468 90244 263474 90256
rect 356698 90244 356704 90256
rect 356756 90244 356762 90296
rect 257890 90176 257896 90228
rect 257948 90216 257954 90228
rect 339494 90216 339500 90228
rect 257948 90188 339500 90216
rect 257948 90176 257954 90188
rect 339494 90176 339500 90188
rect 339552 90176 339558 90228
rect 256326 90108 256332 90160
rect 256384 90148 256390 90160
rect 335354 90148 335360 90160
rect 256384 90120 335360 90148
rect 256384 90108 256390 90120
rect 335354 90108 335360 90120
rect 335412 90108 335418 90160
rect 253566 90040 253572 90092
rect 253624 90080 253630 90092
rect 317414 90080 317420 90092
rect 253624 90052 317420 90080
rect 253624 90040 253630 90052
rect 317414 90040 317420 90052
rect 317472 90040 317478 90092
rect 258994 89632 259000 89684
rect 259052 89672 259058 89684
rect 346394 89672 346400 89684
rect 259052 89644 346400 89672
rect 259052 89632 259058 89644
rect 346394 89632 346400 89644
rect 346452 89632 346458 89684
rect 265986 89564 265992 89616
rect 266044 89604 266050 89616
rect 385678 89604 385684 89616
rect 266044 89576 385684 89604
rect 266044 89564 266050 89576
rect 385678 89564 385684 89576
rect 385736 89564 385742 89616
rect 124122 89496 124128 89548
rect 124180 89536 124186 89548
rect 221274 89536 221280 89548
rect 124180 89508 221280 89536
rect 124180 89496 124186 89508
rect 221274 89496 221280 89508
rect 221332 89496 221338 89548
rect 271690 89496 271696 89548
rect 271748 89536 271754 89548
rect 410518 89536 410524 89548
rect 271748 89508 410524 89536
rect 271748 89496 271754 89508
rect 410518 89496 410524 89508
rect 410576 89496 410582 89548
rect 116578 89428 116584 89480
rect 116636 89468 116642 89480
rect 218514 89468 218520 89480
rect 116636 89440 218520 89468
rect 116636 89428 116642 89440
rect 218514 89428 218520 89440
rect 218572 89428 218578 89480
rect 275646 89428 275652 89480
rect 275704 89468 275710 89480
rect 442258 89468 442264 89480
rect 275704 89440 442264 89468
rect 275704 89428 275710 89440
rect 442258 89428 442264 89440
rect 442316 89428 442322 89480
rect 103422 89360 103428 89412
rect 103480 89400 103486 89412
rect 216858 89400 216864 89412
rect 103480 89372 216864 89400
rect 103480 89360 103486 89372
rect 216858 89360 216864 89372
rect 216916 89360 216922 89412
rect 285306 89360 285312 89412
rect 285364 89400 285370 89412
rect 506474 89400 506480 89412
rect 285364 89372 506480 89400
rect 285364 89360 285370 89372
rect 506474 89360 506480 89372
rect 506532 89360 506538 89412
rect 80698 89292 80704 89344
rect 80756 89332 80762 89344
rect 211706 89332 211712 89344
rect 80756 89304 211712 89332
rect 80756 89292 80762 89304
rect 211706 89292 211712 89304
rect 211764 89292 211770 89344
rect 286778 89292 286784 89344
rect 286836 89332 286842 89344
rect 511258 89332 511264 89344
rect 286836 89304 511264 89332
rect 286836 89292 286842 89304
rect 511258 89292 511264 89304
rect 511316 89292 511322 89344
rect 79318 89224 79324 89276
rect 79376 89264 79382 89276
rect 212994 89264 213000 89276
rect 79376 89236 213000 89264
rect 79376 89224 79382 89236
rect 212994 89224 213000 89236
rect 213052 89224 213058 89276
rect 288066 89224 288072 89276
rect 288124 89264 288130 89276
rect 518158 89264 518164 89276
rect 288124 89236 518164 89264
rect 288124 89224 288130 89236
rect 518158 89224 518164 89236
rect 518216 89224 518222 89276
rect 70210 89156 70216 89208
rect 70268 89196 70274 89208
rect 211522 89196 211528 89208
rect 70268 89168 211528 89196
rect 70268 89156 70274 89168
rect 211522 89156 211528 89168
rect 211580 89156 211586 89208
rect 288250 89156 288256 89208
rect 288308 89196 288314 89208
rect 522298 89196 522304 89208
rect 288308 89168 522304 89196
rect 288308 89156 288314 89168
rect 522298 89156 522304 89168
rect 522356 89156 522362 89208
rect 47578 89088 47584 89140
rect 47636 89128 47642 89140
rect 204714 89128 204720 89140
rect 47636 89100 204720 89128
rect 47636 89088 47642 89100
rect 204714 89088 204720 89100
rect 204772 89088 204778 89140
rect 289446 89088 289452 89140
rect 289504 89128 289510 89140
rect 529198 89128 529204 89140
rect 289504 89100 529204 89128
rect 289504 89088 289510 89100
rect 529198 89088 529204 89100
rect 529256 89088 529262 89140
rect 35158 89020 35164 89072
rect 35216 89060 35222 89072
rect 203150 89060 203156 89072
rect 35216 89032 203156 89060
rect 35216 89020 35222 89032
rect 203150 89020 203156 89032
rect 203208 89020 203214 89072
rect 290918 89020 290924 89072
rect 290976 89060 290982 89072
rect 538214 89060 538220 89072
rect 290976 89032 538220 89060
rect 290976 89020 290982 89032
rect 538214 89020 538220 89032
rect 538272 89020 538278 89072
rect 21358 88952 21364 89004
rect 21416 88992 21422 89004
rect 201770 88992 201776 89004
rect 21416 88964 201776 88992
rect 21416 88952 21422 88964
rect 201770 88952 201776 88964
rect 201828 88952 201834 89004
rect 248138 88952 248144 89004
rect 248196 88992 248202 89004
rect 287054 88992 287060 89004
rect 248196 88964 287060 88992
rect 248196 88952 248202 88964
rect 287054 88952 287060 88964
rect 287112 88952 287118 89004
rect 296346 88952 296352 89004
rect 296404 88992 296410 89004
rect 569954 88992 569960 89004
rect 296404 88964 569960 88992
rect 296404 88952 296410 88964
rect 569954 88952 569960 88964
rect 570012 88952 570018 89004
rect 257706 88884 257712 88936
rect 257764 88924 257770 88936
rect 342254 88924 342260 88936
rect 257764 88896 342260 88924
rect 257764 88884 257770 88896
rect 342254 88884 342260 88896
rect 342312 88884 342318 88936
rect 256418 88816 256424 88868
rect 256476 88856 256482 88868
rect 331858 88856 331864 88868
rect 256476 88828 331864 88856
rect 256476 88816 256482 88828
rect 331858 88816 331864 88828
rect 331916 88816 331922 88868
rect 253658 88748 253664 88800
rect 253716 88788 253722 88800
rect 311250 88788 311256 88800
rect 253716 88760 311256 88788
rect 253716 88748 253722 88760
rect 311250 88748 311256 88760
rect 311308 88748 311314 88800
rect 261938 88272 261944 88324
rect 261996 88312 262002 88324
rect 360194 88312 360200 88324
rect 261996 88284 360200 88312
rect 261996 88272 262002 88284
rect 360194 88272 360200 88284
rect 360252 88272 360258 88324
rect 262030 88204 262036 88256
rect 262088 88244 262094 88256
rect 364334 88244 364340 88256
rect 262088 88216 364340 88244
rect 262088 88204 262094 88216
rect 364334 88204 364340 88216
rect 364392 88204 364398 88256
rect 263502 88136 263508 88188
rect 263560 88176 263566 88188
rect 374086 88176 374092 88188
rect 263560 88148 374092 88176
rect 263560 88136 263566 88148
rect 374086 88136 374092 88148
rect 374144 88136 374150 88188
rect 264698 88068 264704 88120
rect 264756 88108 264762 88120
rect 378134 88108 378140 88120
rect 264756 88080 378140 88108
rect 264756 88068 264762 88080
rect 378134 88068 378140 88080
rect 378192 88068 378198 88120
rect 267182 88000 267188 88052
rect 267240 88040 267246 88052
rect 392578 88040 392584 88052
rect 267240 88012 392584 88040
rect 267240 88000 267246 88012
rect 392578 88000 392584 88012
rect 392636 88000 392642 88052
rect 111058 87932 111064 87984
rect 111116 87972 111122 87984
rect 218330 87972 218336 87984
rect 111116 87944 218336 87972
rect 111116 87932 111122 87944
rect 218330 87932 218336 87944
rect 218388 87932 218394 87984
rect 273070 87932 273076 87984
rect 273128 87972 273134 87984
rect 427814 87972 427820 87984
rect 273128 87944 427820 87972
rect 273128 87932 273134 87944
rect 427814 87932 427820 87944
rect 427872 87932 427878 87984
rect 88978 87864 88984 87916
rect 89036 87904 89042 87916
rect 208946 87904 208952 87916
rect 89036 87876 208952 87904
rect 89036 87864 89042 87876
rect 208946 87864 208952 87876
rect 209004 87864 209010 87916
rect 274174 87864 274180 87916
rect 274232 87904 274238 87916
rect 438854 87904 438860 87916
rect 274232 87876 438860 87904
rect 274232 87864 274238 87876
rect 438854 87864 438860 87876
rect 438912 87864 438918 87916
rect 87598 87796 87604 87848
rect 87656 87836 87662 87848
rect 208578 87836 208584 87848
rect 87656 87808 208584 87836
rect 87656 87796 87662 87808
rect 208578 87796 208584 87808
rect 208636 87796 208642 87848
rect 293678 87796 293684 87848
rect 293736 87836 293742 87848
rect 536098 87836 536104 87848
rect 293736 87808 536104 87836
rect 293736 87796 293742 87808
rect 536098 87796 536104 87808
rect 536156 87796 536162 87848
rect 86218 87728 86224 87780
rect 86276 87768 86282 87780
rect 212902 87768 212908 87780
rect 86276 87740 212908 87768
rect 86276 87728 86282 87740
rect 212902 87728 212908 87740
rect 212960 87728 212966 87780
rect 292298 87728 292304 87780
rect 292356 87768 292362 87780
rect 542998 87768 543004 87780
rect 292356 87740 543004 87768
rect 292356 87728 292362 87740
rect 542998 87728 543004 87740
rect 543056 87728 543062 87780
rect 44082 87660 44088 87712
rect 44140 87700 44146 87712
rect 203518 87700 203524 87712
rect 44140 87672 203524 87700
rect 44140 87660 44146 87672
rect 203518 87660 203524 87672
rect 203576 87660 203582 87712
rect 292206 87660 292212 87712
rect 292264 87700 292270 87712
rect 547966 87700 547972 87712
rect 292264 87672 547972 87700
rect 292264 87660 292270 87672
rect 547966 87660 547972 87672
rect 548024 87660 548030 87712
rect 15838 87592 15844 87644
rect 15896 87632 15902 87644
rect 202322 87632 202328 87644
rect 15896 87604 202328 87632
rect 15896 87592 15902 87604
rect 202322 87592 202328 87604
rect 202380 87592 202386 87644
rect 296438 87592 296444 87644
rect 296496 87632 296502 87644
rect 565814 87632 565820 87644
rect 296496 87604 565820 87632
rect 296496 87592 296502 87604
rect 565814 87592 565820 87604
rect 565872 87592 565878 87644
rect 260466 87524 260472 87576
rect 260524 87564 260530 87576
rect 357434 87564 357440 87576
rect 260524 87536 357440 87564
rect 260524 87524 260530 87536
rect 357434 87524 357440 87536
rect 357492 87524 357498 87576
rect 311158 86912 311164 86964
rect 311216 86952 311222 86964
rect 580166 86952 580172 86964
rect 311216 86924 580172 86952
rect 311216 86912 311222 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 261754 86844 261760 86896
rect 261812 86884 261818 86896
rect 367094 86884 367100 86896
rect 261812 86856 367100 86884
rect 261812 86844 261818 86856
rect 367094 86844 367100 86856
rect 367152 86844 367158 86896
rect 270034 86776 270040 86828
rect 270092 86816 270098 86828
rect 381538 86816 381544 86828
rect 270092 86788 381544 86816
rect 270092 86776 270098 86788
rect 381538 86776 381544 86788
rect 381596 86776 381602 86828
rect 264422 86708 264428 86760
rect 264480 86748 264486 86760
rect 382366 86748 382372 86760
rect 264480 86720 382372 86748
rect 264480 86708 264486 86720
rect 382366 86708 382372 86720
rect 382424 86708 382430 86760
rect 267274 86640 267280 86692
rect 267332 86680 267338 86692
rect 395338 86680 395344 86692
rect 267332 86652 395344 86680
rect 267332 86640 267338 86652
rect 395338 86640 395344 86652
rect 395396 86640 395402 86692
rect 272794 86572 272800 86624
rect 272852 86612 272858 86624
rect 406378 86612 406384 86624
rect 272852 86584 406384 86612
rect 272852 86572 272858 86584
rect 406378 86572 406384 86584
rect 406436 86572 406442 86624
rect 274266 86504 274272 86556
rect 274324 86544 274330 86556
rect 441614 86544 441620 86556
rect 274324 86516 441620 86544
rect 274324 86504 274330 86516
rect 441614 86504 441620 86516
rect 441672 86504 441678 86556
rect 122098 86436 122104 86488
rect 122156 86476 122162 86488
rect 217410 86476 217416 86488
rect 122156 86448 217416 86476
rect 122156 86436 122162 86448
rect 217410 86436 217416 86448
rect 217468 86436 217474 86488
rect 275738 86436 275744 86488
rect 275796 86476 275802 86488
rect 448606 86476 448612 86488
rect 275796 86448 448612 86476
rect 275796 86436 275802 86448
rect 448606 86436 448612 86448
rect 448664 86436 448670 86488
rect 33042 86368 33048 86420
rect 33100 86408 33106 86420
rect 199378 86408 199384 86420
rect 33100 86380 199384 86408
rect 33100 86368 33106 86380
rect 199378 86368 199384 86380
rect 199436 86368 199442 86420
rect 279970 86368 279976 86420
rect 280028 86408 280034 86420
rect 470594 86408 470600 86420
rect 280028 86380 470600 86408
rect 280028 86368 280034 86380
rect 470594 86368 470600 86380
rect 470652 86368 470658 86420
rect 28258 86300 28264 86352
rect 28316 86340 28322 86352
rect 201586 86340 201592 86352
rect 28316 86312 201592 86340
rect 28316 86300 28322 86312
rect 201586 86300 201592 86312
rect 201644 86300 201650 86352
rect 284110 86300 284116 86352
rect 284168 86340 284174 86352
rect 496814 86340 496820 86352
rect 284168 86312 496820 86340
rect 284168 86300 284174 86312
rect 496814 86300 496820 86312
rect 496872 86300 496878 86352
rect 5442 86232 5448 86284
rect 5500 86272 5506 86284
rect 195330 86272 195336 86284
rect 5500 86244 195336 86272
rect 5500 86232 5506 86244
rect 195330 86232 195336 86244
rect 195388 86232 195394 86284
rect 290458 86232 290464 86284
rect 290516 86272 290522 86284
rect 535454 86272 535460 86284
rect 290516 86244 535460 86272
rect 290516 86232 290522 86244
rect 535454 86232 535460 86244
rect 535512 86232 535518 86284
rect 256142 86164 256148 86216
rect 256200 86204 256206 86216
rect 329834 86204 329840 86216
rect 256200 86176 329840 86204
rect 256200 86164 256206 86176
rect 329834 86164 329840 86176
rect 329892 86164 329898 86216
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 151078 85524 151084 85536
rect 3200 85496 151084 85524
rect 3200 85484 3206 85496
rect 151078 85484 151084 85496
rect 151136 85484 151142 85536
rect 253382 85416 253388 85468
rect 253440 85456 253446 85468
rect 318058 85456 318064 85468
rect 253440 85428 318064 85456
rect 253440 85416 253446 85428
rect 318058 85416 318064 85428
rect 318116 85416 318122 85468
rect 263042 85348 263048 85400
rect 263100 85388 263106 85400
rect 340966 85388 340972 85400
rect 263100 85360 340972 85388
rect 263100 85348 263106 85360
rect 340966 85348 340972 85360
rect 341024 85348 341030 85400
rect 259086 85280 259092 85332
rect 259144 85320 259150 85332
rect 342898 85320 342904 85332
rect 259144 85292 342904 85320
rect 259144 85280 259150 85292
rect 342898 85280 342904 85292
rect 342956 85280 342962 85332
rect 271322 85212 271328 85264
rect 271380 85252 271386 85264
rect 375374 85252 375380 85264
rect 271380 85224 375380 85252
rect 271380 85212 271386 85224
rect 375374 85212 375380 85224
rect 375432 85212 375438 85264
rect 279786 85144 279792 85196
rect 279844 85184 279850 85196
rect 472710 85184 472716 85196
rect 279844 85156 472716 85184
rect 279844 85144 279850 85156
rect 472710 85144 472716 85156
rect 472768 85144 472774 85196
rect 281902 85076 281908 85128
rect 281960 85116 281966 85128
rect 482278 85116 482284 85128
rect 281960 85088 482284 85116
rect 281960 85076 281966 85088
rect 482278 85076 482284 85088
rect 482336 85076 482342 85128
rect 283834 85008 283840 85060
rect 283892 85048 283898 85060
rect 492674 85048 492680 85060
rect 283892 85020 492680 85048
rect 283892 85008 283898 85020
rect 492674 85008 492680 85020
rect 492732 85008 492738 85060
rect 285490 84940 285496 84992
rect 285548 84980 285554 84992
rect 499574 84980 499580 84992
rect 285548 84952 499580 84980
rect 285548 84940 285554 84952
rect 499574 84940 499580 84952
rect 499632 84940 499638 84992
rect 289538 84872 289544 84924
rect 289596 84912 289602 84924
rect 524414 84912 524420 84924
rect 289596 84884 524420 84912
rect 289596 84872 289602 84884
rect 524414 84872 524420 84884
rect 524472 84872 524478 84924
rect 107562 84804 107568 84856
rect 107620 84844 107626 84856
rect 196618 84844 196624 84856
rect 107620 84816 196624 84844
rect 107620 84804 107626 84816
rect 196618 84804 196624 84816
rect 196676 84804 196682 84856
rect 293770 84804 293776 84856
rect 293828 84844 293834 84856
rect 553394 84844 553400 84856
rect 293828 84816 553400 84844
rect 293828 84804 293834 84816
rect 553394 84804 553400 84816
rect 553452 84804 553458 84856
rect 276658 83852 276664 83904
rect 276716 83892 276722 83904
rect 357526 83892 357532 83904
rect 276716 83864 357532 83892
rect 276716 83852 276722 83864
rect 357526 83852 357532 83864
rect 357584 83852 357590 83904
rect 262950 83784 262956 83836
rect 263008 83824 263014 83836
rect 365806 83824 365812 83836
rect 263008 83796 365812 83824
rect 263008 83784 263014 83796
rect 365806 83784 365812 83796
rect 365864 83784 365870 83836
rect 274358 83716 274364 83768
rect 274416 83756 274422 83768
rect 418798 83756 418804 83768
rect 274416 83728 418804 83756
rect 274416 83716 274422 83728
rect 418798 83716 418804 83728
rect 418856 83716 418862 83768
rect 286502 83648 286508 83700
rect 286560 83688 286566 83700
rect 510614 83688 510620 83700
rect 286560 83660 510620 83688
rect 286560 83648 286566 83660
rect 510614 83648 510620 83660
rect 510672 83648 510678 83700
rect 287882 83580 287888 83632
rect 287940 83620 287946 83632
rect 517514 83620 517520 83632
rect 287940 83592 517520 83620
rect 287940 83580 287946 83592
rect 517514 83580 517520 83592
rect 517572 83580 517578 83632
rect 290826 83512 290832 83564
rect 290884 83552 290890 83564
rect 539686 83552 539692 83564
rect 290884 83524 539692 83552
rect 290884 83512 290890 83524
rect 539686 83512 539692 83524
rect 539744 83512 539750 83564
rect 246666 83444 246672 83496
rect 246724 83484 246730 83496
rect 273898 83484 273904 83496
rect 246724 83456 273904 83484
rect 246724 83444 246730 83456
rect 273898 83444 273904 83456
rect 273956 83444 273962 83496
rect 293586 83444 293592 83496
rect 293644 83484 293650 83496
rect 556246 83484 556252 83496
rect 293644 83456 556252 83484
rect 293644 83444 293650 83456
rect 556246 83444 556252 83456
rect 556304 83444 556310 83496
rect 298830 82424 298836 82476
rect 298888 82464 298894 82476
rect 400214 82464 400220 82476
rect 298888 82436 400220 82464
rect 298888 82424 298894 82436
rect 400214 82424 400220 82436
rect 400272 82424 400278 82476
rect 264514 82356 264520 82408
rect 264572 82396 264578 82408
rect 377398 82396 377404 82408
rect 264572 82368 377404 82396
rect 264572 82356 264578 82368
rect 377398 82356 377404 82368
rect 377456 82356 377462 82408
rect 275830 82288 275836 82340
rect 275888 82328 275894 82340
rect 396718 82328 396724 82340
rect 275888 82300 396724 82328
rect 275888 82288 275894 82300
rect 396718 82288 396724 82300
rect 396776 82288 396782 82340
rect 271782 82220 271788 82272
rect 271840 82260 271846 82272
rect 393958 82260 393964 82272
rect 271840 82232 393964 82260
rect 271840 82220 271846 82232
rect 393958 82220 393964 82232
rect 394016 82220 394022 82272
rect 296162 82152 296168 82204
rect 296220 82192 296226 82204
rect 565078 82192 565084 82204
rect 296220 82164 565084 82192
rect 296220 82152 296226 82164
rect 565078 82152 565084 82164
rect 565136 82152 565142 82204
rect 248230 82084 248236 82136
rect 248288 82124 248294 82136
rect 275278 82124 275284 82136
rect 248288 82096 275284 82124
rect 248288 82084 248294 82096
rect 275278 82084 275284 82096
rect 275336 82084 275342 82136
rect 278498 82084 278504 82136
rect 278556 82124 278562 82136
rect 295978 82124 295984 82136
rect 278556 82096 295984 82124
rect 278556 82084 278562 82096
rect 295978 82084 295984 82096
rect 296036 82084 296042 82136
rect 304350 82084 304356 82136
rect 304408 82124 304414 82136
rect 582558 82124 582564 82136
rect 304408 82096 582564 82124
rect 304408 82084 304414 82096
rect 582558 82084 582564 82096
rect 582616 82084 582622 82136
rect 275554 80792 275560 80844
rect 275612 80832 275618 80844
rect 399478 80832 399484 80844
rect 275612 80804 399484 80832
rect 275612 80792 275618 80804
rect 399478 80792 399484 80804
rect 399536 80792 399542 80844
rect 274450 80724 274456 80776
rect 274508 80764 274514 80776
rect 411898 80764 411904 80776
rect 274508 80736 411904 80764
rect 274508 80724 274514 80736
rect 411898 80724 411904 80736
rect 411956 80724 411962 80776
rect 248046 80656 248052 80708
rect 248104 80696 248110 80708
rect 284294 80696 284300 80708
rect 248104 80668 284300 80696
rect 248104 80656 248110 80668
rect 284294 80656 284300 80668
rect 284352 80656 284358 80708
rect 298738 80656 298744 80708
rect 298796 80696 298802 80708
rect 575474 80696 575480 80708
rect 298796 80668 575480 80696
rect 298796 80656 298802 80668
rect 575474 80656 575480 80668
rect 575532 80656 575538 80708
rect 316678 73108 316684 73160
rect 316736 73148 316742 73160
rect 579982 73148 579988 73160
rect 316736 73120 579988 73148
rect 316736 73108 316742 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 253474 72428 253480 72480
rect 253532 72468 253538 72480
rect 316126 72468 316132 72480
rect 253532 72440 316132 72468
rect 253532 72428 253538 72440
rect 316126 72428 316132 72440
rect 316184 72428 316190 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 157978 71720 157984 71732
rect 3476 71692 157984 71720
rect 3476 71680 3482 71692
rect 157978 71680 157984 71692
rect 158036 71680 158042 71732
rect 530578 60664 530584 60716
rect 530636 60704 530642 60716
rect 580166 60704 580172 60716
rect 530636 60676 580172 60704
rect 530636 60664 530642 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 289170 59984 289176 60036
rect 289228 60024 289234 60036
rect 530670 60024 530676 60036
rect 289228 59996 530676 60024
rect 289228 59984 289234 59996
rect 530670 59984 530676 59996
rect 530728 59984 530734 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 32398 59344 32404 59356
rect 3108 59316 32404 59344
rect 3108 59304 3114 59316
rect 32398 59304 32404 59316
rect 32456 59304 32462 59356
rect 68922 47540 68928 47592
rect 68980 47580 68986 47592
rect 197998 47580 198004 47592
rect 68980 47552 198004 47580
rect 68980 47540 68986 47552
rect 197998 47540 198004 47552
rect 198056 47540 198062 47592
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 148318 45540 148324 45552
rect 3476 45512 148324 45540
rect 3476 45500 3482 45512
rect 148318 45500 148324 45512
rect 148376 45500 148382 45552
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 156598 33096 156604 33108
rect 3200 33068 156604 33096
rect 3200 33056 3206 33068
rect 156598 33056 156604 33068
rect 156656 33056 156662 33108
rect 313918 33056 313924 33108
rect 313976 33096 313982 33108
rect 580166 33096 580172 33108
rect 313976 33068 580172 33096
rect 313976 33056 313982 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 286594 26868 286600 26920
rect 286652 26908 286658 26920
rect 514846 26908 514852 26920
rect 286652 26880 514852 26908
rect 286652 26868 286658 26880
rect 514846 26868 514852 26880
rect 514904 26868 514910 26920
rect 285030 24080 285036 24132
rect 285088 24120 285094 24132
rect 506566 24120 506572 24132
rect 285088 24092 506572 24120
rect 285088 24080 285094 24092
rect 506566 24080 506572 24092
rect 506624 24080 506630 24132
rect 296254 22720 296260 22772
rect 296312 22760 296318 22772
rect 571334 22760 571340 22772
rect 296312 22732 571340 22760
rect 296312 22720 296318 22732
rect 571334 22720 571340 22732
rect 571392 22720 571398 22772
rect 292022 21360 292028 21412
rect 292080 21400 292086 21412
rect 546494 21400 546500 21412
rect 292080 21372 546500 21400
rect 292080 21360 292086 21372
rect 546494 21360 546500 21372
rect 546552 21360 546558 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 43438 20652 43444 20664
rect 3476 20624 43444 20652
rect 3476 20612 3482 20624
rect 43438 20612 43444 20624
rect 43496 20612 43502 20664
rect 525058 20612 525064 20664
rect 525116 20652 525122 20664
rect 580166 20652 580172 20664
rect 525116 20624 580172 20652
rect 525116 20612 525122 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 282454 19932 282460 19984
rect 282512 19972 282518 19984
rect 490006 19972 490012 19984
rect 282512 19944 490012 19972
rect 282512 19932 282518 19944
rect 490006 19932 490012 19944
rect 490064 19932 490070 19984
rect 188982 18572 188988 18624
rect 189040 18612 189046 18624
rect 230842 18612 230848 18624
rect 189040 18584 230848 18612
rect 189040 18572 189046 18584
rect 230842 18572 230848 18584
rect 230900 18572 230906 18624
rect 287974 18572 287980 18624
rect 288032 18612 288038 18624
rect 521654 18612 521660 18624
rect 288032 18584 521660 18612
rect 288032 18572 288038 18584
rect 521654 18572 521660 18584
rect 521712 18572 521718 18624
rect 250806 16056 250812 16108
rect 250864 16096 250870 16108
rect 298094 16096 298100 16108
rect 250864 16068 298100 16096
rect 250864 16056 250870 16068
rect 298094 16056 298100 16068
rect 298152 16056 298158 16108
rect 250898 15988 250904 16040
rect 250956 16028 250962 16040
rect 301498 16028 301504 16040
rect 250956 16000 301504 16028
rect 250956 15988 250962 16000
rect 301498 15988 301504 16000
rect 301556 15988 301562 16040
rect 252094 15920 252100 15972
rect 252152 15960 252158 15972
rect 307754 15960 307760 15972
rect 252152 15932 307760 15960
rect 252152 15920 252158 15932
rect 307754 15920 307760 15932
rect 307812 15920 307818 15972
rect 106182 15852 106188 15904
rect 106240 15892 106246 15904
rect 217134 15892 217140 15904
rect 106240 15864 217140 15892
rect 106240 15852 106246 15864
rect 217134 15852 217140 15864
rect 217192 15852 217198 15904
rect 240042 15852 240048 15904
rect 240100 15892 240106 15904
rect 253474 15892 253480 15904
rect 240100 15864 253480 15892
rect 240100 15852 240106 15864
rect 253474 15852 253480 15864
rect 253532 15852 253538 15904
rect 254854 15852 254860 15904
rect 254912 15892 254918 15904
rect 322934 15892 322940 15904
rect 254912 15864 322940 15892
rect 254912 15852 254918 15864
rect 322934 15852 322940 15864
rect 322992 15852 322998 15904
rect 323578 15852 323584 15904
rect 323636 15892 323642 15904
rect 404354 15892 404360 15904
rect 323636 15864 404360 15892
rect 323636 15852 323642 15864
rect 404354 15852 404360 15864
rect 404412 15852 404418 15904
rect 294966 14628 294972 14680
rect 295024 14668 295030 14680
rect 560386 14668 560392 14680
rect 295024 14640 560392 14668
rect 295024 14628 295030 14640
rect 560386 14628 560392 14640
rect 560444 14628 560450 14680
rect 294874 14560 294880 14612
rect 294932 14600 294938 14612
rect 564434 14600 564440 14612
rect 294932 14572 564440 14600
rect 294932 14560 294938 14572
rect 564434 14560 564440 14572
rect 564492 14560 564498 14612
rect 297818 14492 297824 14544
rect 297876 14532 297882 14544
rect 575106 14532 575112 14544
rect 297876 14504 575112 14532
rect 297876 14492 297882 14504
rect 575106 14492 575112 14504
rect 575164 14492 575170 14544
rect 161198 14424 161204 14476
rect 161256 14464 161262 14476
rect 226610 14464 226616 14476
rect 161256 14436 226616 14464
rect 161256 14424 161262 14436
rect 226610 14424 226616 14436
rect 226668 14424 226674 14476
rect 258718 14424 258724 14476
rect 258776 14464 258782 14476
rect 281534 14464 281540 14476
rect 258776 14436 281540 14464
rect 258776 14424 258782 14436
rect 281534 14424 281540 14436
rect 281592 14424 281598 14476
rect 297726 14424 297732 14476
rect 297784 14464 297790 14476
rect 578602 14464 578608 14476
rect 297784 14436 578608 14464
rect 297784 14424 297790 14436
rect 578602 14424 578608 14436
rect 578660 14424 578666 14476
rect 256234 13472 256240 13524
rect 256292 13512 256298 13524
rect 333882 13512 333888 13524
rect 256292 13484 333888 13512
rect 256292 13472 256298 13484
rect 333882 13472 333888 13484
rect 333940 13472 333946 13524
rect 277210 13404 277216 13456
rect 277268 13444 277274 13456
rect 453206 13444 453212 13456
rect 277268 13416 453212 13444
rect 277268 13404 277274 13416
rect 453206 13404 453212 13416
rect 453264 13404 453270 13456
rect 277118 13336 277124 13388
rect 277176 13376 277182 13388
rect 456886 13376 456892 13388
rect 277176 13348 456892 13376
rect 277176 13336 277182 13348
rect 456886 13336 456892 13348
rect 456944 13336 456950 13388
rect 278590 13268 278596 13320
rect 278648 13308 278654 13320
rect 459922 13308 459928 13320
rect 278648 13280 459928 13308
rect 278648 13268 278654 13280
rect 459922 13268 459928 13280
rect 459980 13268 459986 13320
rect 278314 13200 278320 13252
rect 278372 13240 278378 13252
rect 463970 13240 463976 13252
rect 278372 13212 463976 13240
rect 278372 13200 278378 13212
rect 463970 13200 463976 13212
rect 464028 13200 464034 13252
rect 281166 13132 281172 13184
rect 281224 13172 281230 13184
rect 478138 13172 478144 13184
rect 281224 13144 478144 13172
rect 281224 13132 281230 13144
rect 478138 13132 478144 13144
rect 478196 13132 478202 13184
rect 170766 13064 170772 13116
rect 170824 13104 170830 13116
rect 228082 13104 228088 13116
rect 170824 13076 228088 13104
rect 170824 13064 170830 13076
rect 228082 13064 228088 13076
rect 228140 13064 228146 13116
rect 246758 13064 246764 13116
rect 246816 13104 246822 13116
rect 266998 13104 267004 13116
rect 246816 13076 267004 13104
rect 246816 13064 246822 13076
rect 266998 13064 267004 13076
rect 267056 13064 267062 13116
rect 281074 13064 281080 13116
rect 281132 13104 281138 13116
rect 482186 13104 482192 13116
rect 281132 13076 482192 13104
rect 281132 13064 281138 13076
rect 482186 13064 482192 13076
rect 482244 13064 482250 13116
rect 266078 12248 266084 12300
rect 266136 12288 266142 12300
rect 385586 12288 385592 12300
rect 266136 12260 385592 12288
rect 266136 12248 266142 12260
rect 385586 12248 385592 12260
rect 385644 12248 385650 12300
rect 266170 12180 266176 12232
rect 266228 12220 266234 12232
rect 389450 12220 389456 12232
rect 266228 12192 389456 12220
rect 266228 12180 266234 12192
rect 389450 12180 389456 12192
rect 389508 12180 389514 12232
rect 265894 12112 265900 12164
rect 265952 12152 265958 12164
rect 392578 12152 392584 12164
rect 265952 12124 392584 12152
rect 265952 12112 265958 12124
rect 392578 12112 392584 12124
rect 392636 12112 392642 12164
rect 267366 12044 267372 12096
rect 267424 12084 267430 12096
rect 396074 12084 396080 12096
rect 267424 12056 396080 12084
rect 267424 12044 267430 12056
rect 396074 12044 396080 12056
rect 396132 12044 396138 12096
rect 267458 11976 267464 12028
rect 267516 12016 267522 12028
rect 398834 12016 398840 12028
rect 267516 11988 398840 12016
rect 267516 11976 267522 11988
rect 398834 11976 398840 11988
rect 398892 11976 398898 12028
rect 268654 11908 268660 11960
rect 268712 11948 268718 11960
rect 403526 11948 403532 11960
rect 268712 11920 403532 11948
rect 268712 11908 268718 11920
rect 403526 11908 403532 11920
rect 403584 11908 403590 11960
rect 268746 11840 268752 11892
rect 268804 11880 268810 11892
rect 407206 11880 407212 11892
rect 268804 11852 407212 11880
rect 268804 11840 268810 11852
rect 407206 11840 407212 11852
rect 407264 11840 407270 11892
rect 245194 11772 245200 11824
rect 245252 11812 245258 11824
rect 256050 11812 256056 11824
rect 245252 11784 256056 11812
rect 245252 11772 245258 11784
rect 256050 11772 256056 11784
rect 256108 11772 256114 11824
rect 270126 11772 270132 11824
rect 270184 11812 270190 11824
rect 410426 11812 410432 11824
rect 270184 11784 410432 11812
rect 270184 11772 270190 11784
rect 410426 11772 410432 11784
rect 410484 11772 410490 11824
rect 111702 11704 111708 11756
rect 111760 11744 111766 11756
rect 119338 11744 119344 11756
rect 111760 11716 119344 11744
rect 111760 11704 111766 11716
rect 119338 11704 119344 11716
rect 119396 11704 119402 11756
rect 119890 11704 119896 11756
rect 119948 11744 119954 11756
rect 219894 11744 219900 11756
rect 119948 11716 219900 11744
rect 119948 11704 119954 11716
rect 219894 11704 219900 11716
rect 219952 11704 219958 11756
rect 243906 11704 243912 11756
rect 243964 11744 243970 11756
rect 256142 11744 256148 11756
rect 243964 11716 256148 11744
rect 243964 11704 243970 11716
rect 256142 11704 256148 11716
rect 256200 11704 256206 11756
rect 270218 11704 270224 11756
rect 270276 11744 270282 11756
rect 414290 11744 414296 11756
rect 270276 11716 414296 11744
rect 270276 11704 270282 11716
rect 414290 11704 414296 11716
rect 414348 11704 414354 11756
rect 357526 11636 357532 11688
rect 357584 11676 357590 11688
rect 358722 11676 358728 11688
rect 357584 11648 358728 11676
rect 357584 11636 357590 11648
rect 358722 11636 358728 11648
rect 358780 11636 358786 11688
rect 250990 10888 250996 10940
rect 251048 10928 251054 10940
rect 299566 10928 299572 10940
rect 251048 10900 299572 10928
rect 251048 10888 251054 10900
rect 299566 10888 299572 10900
rect 299624 10888 299630 10940
rect 252186 10820 252192 10872
rect 252244 10860 252250 10872
rect 303890 10860 303896 10872
rect 252244 10832 303896 10860
rect 252244 10820 252250 10832
rect 303890 10820 303896 10832
rect 303948 10820 303954 10872
rect 252278 10752 252284 10804
rect 252336 10792 252342 10804
rect 307938 10792 307944 10804
rect 252336 10764 307944 10792
rect 252336 10752 252342 10764
rect 307938 10752 307944 10764
rect 307996 10752 308002 10804
rect 252370 10684 252376 10736
rect 252428 10724 252434 10736
rect 311158 10724 311164 10736
rect 252428 10696 311164 10724
rect 252428 10684 252434 10696
rect 311158 10684 311164 10696
rect 311216 10684 311222 10736
rect 117222 10616 117228 10668
rect 117280 10656 117286 10668
rect 220262 10656 220268 10668
rect 117280 10628 220268 10656
rect 117280 10616 117286 10628
rect 220262 10616 220268 10628
rect 220320 10616 220326 10668
rect 255038 10616 255044 10668
rect 255096 10656 255102 10668
rect 322106 10656 322112 10668
rect 255096 10628 322112 10656
rect 255096 10616 255102 10628
rect 322106 10616 322112 10628
rect 322164 10616 322170 10668
rect 99282 10548 99288 10600
rect 99340 10588 99346 10600
rect 215478 10588 215484 10600
rect 99340 10560 215484 10588
rect 99340 10548 99346 10560
rect 215478 10548 215484 10560
rect 215536 10548 215542 10600
rect 254946 10548 254952 10600
rect 255004 10588 255010 10600
rect 324314 10588 324320 10600
rect 255004 10560 324320 10588
rect 255004 10548 255010 10560
rect 324314 10548 324320 10560
rect 324372 10548 324378 10600
rect 95142 10480 95148 10532
rect 95200 10520 95206 10532
rect 216030 10520 216036 10532
rect 95200 10492 216036 10520
rect 95200 10480 95206 10492
rect 216030 10480 216036 10492
rect 216088 10480 216094 10532
rect 295150 10480 295156 10532
rect 295208 10520 295214 10532
rect 559282 10520 559288 10532
rect 295208 10492 559288 10520
rect 295208 10480 295214 10492
rect 559282 10480 559288 10492
rect 559340 10480 559346 10532
rect 92382 10412 92388 10464
rect 92440 10452 92446 10464
rect 215662 10452 215668 10464
rect 92440 10424 215668 10452
rect 92440 10412 92446 10424
rect 215662 10412 215668 10424
rect 215720 10412 215726 10464
rect 295058 10412 295064 10464
rect 295116 10452 295122 10464
rect 563238 10452 563244 10464
rect 295116 10424 563244 10452
rect 295116 10412 295122 10424
rect 563238 10412 563244 10424
rect 563296 10412 563302 10464
rect 87966 10344 87972 10396
rect 88024 10384 88030 10396
rect 214098 10384 214104 10396
rect 88024 10356 214104 10384
rect 88024 10344 88030 10356
rect 214098 10344 214104 10356
rect 214156 10344 214162 10396
rect 298002 10344 298008 10396
rect 298060 10384 298066 10396
rect 573450 10384 573456 10396
rect 298060 10356 573456 10384
rect 298060 10344 298066 10356
rect 573450 10344 573456 10356
rect 573508 10344 573514 10396
rect 85482 10276 85488 10328
rect 85540 10316 85546 10328
rect 214190 10316 214196 10328
rect 85540 10288 214196 10316
rect 85540 10276 85546 10288
rect 214190 10276 214196 10288
rect 214248 10276 214254 10328
rect 297910 10276 297916 10328
rect 297968 10316 297974 10328
rect 576946 10316 576952 10328
rect 297968 10288 576952 10316
rect 297968 10276 297974 10288
rect 576946 10276 576952 10288
rect 577004 10276 577010 10328
rect 122282 9460 122288 9512
rect 122340 9500 122346 9512
rect 219710 9500 219716 9512
rect 122340 9472 219716 9500
rect 122340 9460 122346 9472
rect 219710 9460 219716 9472
rect 219768 9460 219774 9512
rect 118786 9392 118792 9444
rect 118844 9432 118850 9444
rect 219526 9432 219532 9444
rect 118844 9404 219532 9432
rect 118844 9392 118850 9404
rect 219526 9392 219532 9404
rect 219584 9392 219590 9444
rect 115290 9324 115296 9376
rect 115348 9364 115354 9376
rect 220446 9364 220452 9376
rect 115348 9336 220452 9364
rect 115348 9324 115354 9336
rect 220446 9324 220452 9336
rect 220504 9324 220510 9376
rect 97442 9256 97448 9308
rect 97500 9296 97506 9308
rect 215754 9296 215760 9308
rect 97500 9268 215760 9296
rect 97500 9256 97506 9268
rect 215754 9256 215760 9268
rect 215812 9256 215818 9308
rect 93946 9188 93952 9240
rect 94004 9228 94010 9240
rect 215846 9228 215852 9240
rect 94004 9200 215852 9228
rect 94004 9188 94010 9200
rect 215846 9188 215852 9200
rect 215904 9188 215910 9240
rect 90450 9120 90456 9172
rect 90508 9160 90514 9172
rect 214466 9160 214472 9172
rect 90508 9132 214472 9160
rect 90508 9120 90514 9132
rect 214466 9120 214472 9132
rect 214524 9120 214530 9172
rect 86862 9052 86868 9104
rect 86920 9092 86926 9104
rect 214282 9092 214288 9104
rect 86920 9064 214288 9092
rect 86920 9052 86926 9064
rect 214282 9052 214288 9064
rect 214340 9052 214346 9104
rect 300118 9052 300124 9104
rect 300176 9092 300182 9104
rect 362310 9092 362316 9104
rect 300176 9064 362316 9092
rect 300176 9052 300182 9064
rect 362310 9052 362316 9064
rect 362368 9052 362374 9104
rect 33594 8984 33600 9036
rect 33652 9024 33658 9036
rect 205634 9024 205640 9036
rect 33652 8996 205640 9024
rect 33652 8984 33658 8996
rect 205634 8984 205640 8996
rect 205692 8984 205698 9036
rect 281258 8984 281264 9036
rect 281316 9024 281322 9036
rect 476942 9024 476948 9036
rect 281316 8996 476948 9024
rect 281316 8984 281322 8996
rect 476942 8984 476948 8996
rect 477000 8984 477006 9036
rect 30098 8916 30104 8968
rect 30156 8956 30162 8968
rect 204990 8956 204996 8968
rect 30156 8928 204996 8956
rect 30156 8916 30162 8928
rect 204990 8916 204996 8928
rect 205048 8916 205054 8968
rect 220446 8916 220452 8968
rect 220504 8956 220510 8968
rect 231302 8956 231308 8968
rect 220504 8928 231308 8956
rect 220504 8916 220510 8928
rect 231302 8916 231308 8928
rect 231360 8916 231366 8968
rect 253198 8916 253204 8968
rect 253256 8956 253262 8968
rect 280706 8956 280712 8968
rect 253256 8928 280712 8956
rect 253256 8916 253262 8928
rect 280706 8916 280712 8928
rect 280764 8916 280770 8968
rect 281350 8916 281356 8968
rect 281408 8956 281414 8968
rect 481726 8956 481732 8968
rect 281408 8928 481732 8956
rect 281408 8916 281414 8928
rect 481726 8916 481732 8928
rect 481784 8916 481790 8968
rect 260098 8236 260104 8288
rect 260156 8276 260162 8288
rect 264146 8276 264152 8288
rect 260156 8248 264152 8276
rect 260156 8236 260162 8248
rect 264146 8236 264152 8248
rect 264204 8236 264210 8288
rect 202690 8100 202696 8152
rect 202748 8140 202754 8152
rect 233418 8140 233424 8152
rect 202748 8112 233424 8140
rect 202748 8100 202754 8112
rect 233418 8100 233424 8112
rect 233476 8100 233482 8152
rect 199102 8032 199108 8084
rect 199160 8072 199166 8084
rect 233786 8072 233792 8084
rect 199160 8044 233792 8072
rect 199160 8032 199166 8044
rect 233786 8032 233792 8044
rect 233844 8032 233850 8084
rect 267642 8032 267648 8084
rect 267700 8072 267706 8084
rect 395246 8072 395252 8084
rect 267700 8044 395252 8072
rect 267700 8032 267706 8044
rect 395246 8032 395252 8044
rect 395304 8032 395310 8084
rect 142798 8004 142804 8016
rect 142126 7976 142804 8004
rect 74994 7896 75000 7948
rect 75052 7936 75058 7948
rect 142126 7936 142154 7976
rect 142798 7964 142804 7976
rect 142856 7964 142862 8016
rect 195606 7964 195612 8016
rect 195664 8004 195670 8016
rect 232682 8004 232688 8016
rect 195664 7976 232688 8004
rect 195664 7964 195670 7976
rect 232682 7964 232688 7976
rect 232740 7964 232746 8016
rect 267550 7964 267556 8016
rect 267608 8004 267614 8016
rect 398926 8004 398932 8016
rect 267608 7976 398932 8004
rect 267608 7964 267614 7976
rect 398926 7964 398932 7976
rect 398984 7964 398990 8016
rect 75052 7908 142154 7936
rect 75052 7896 75058 7908
rect 142430 7896 142436 7948
rect 142488 7936 142494 7948
rect 223942 7936 223948 7948
rect 142488 7908 223948 7936
rect 142488 7896 142494 7908
rect 223942 7896 223948 7908
rect 224000 7896 224006 7948
rect 268562 7896 268568 7948
rect 268620 7936 268626 7948
rect 402514 7936 402520 7948
rect 268620 7908 402520 7936
rect 268620 7896 268626 7908
rect 402514 7896 402520 7908
rect 402572 7896 402578 7948
rect 222470 7868 222476 7880
rect 142126 7840 222476 7868
rect 138842 7760 138848 7812
rect 138900 7800 138906 7812
rect 142126 7800 142154 7840
rect 222470 7828 222476 7840
rect 222528 7828 222534 7880
rect 268930 7828 268936 7880
rect 268988 7868 268994 7880
rect 406010 7868 406016 7880
rect 268988 7840 406016 7868
rect 268988 7828 268994 7840
rect 406010 7828 406016 7840
rect 406068 7828 406074 7880
rect 138900 7772 142154 7800
rect 138900 7760 138906 7772
rect 146938 7760 146944 7812
rect 146996 7800 147002 7812
rect 222746 7800 222752 7812
rect 146996 7772 222752 7800
rect 146996 7760 147002 7772
rect 222746 7760 222752 7772
rect 222804 7760 222810 7812
rect 268838 7760 268844 7812
rect 268896 7800 268902 7812
rect 409598 7800 409604 7812
rect 268896 7772 409604 7800
rect 268896 7760 268902 7772
rect 409598 7760 409604 7772
rect 409656 7760 409662 7812
rect 131758 7692 131764 7744
rect 131816 7732 131822 7744
rect 222930 7732 222936 7744
rect 131816 7704 222936 7732
rect 131816 7692 131822 7704
rect 222930 7692 222936 7704
rect 222988 7692 222994 7744
rect 270310 7692 270316 7744
rect 270368 7732 270374 7744
rect 413094 7732 413100 7744
rect 270368 7704 413100 7732
rect 270368 7692 270374 7704
rect 413094 7692 413100 7704
rect 413152 7692 413158 7744
rect 50154 7624 50160 7676
rect 50212 7664 50218 7676
rect 192478 7664 192484 7676
rect 50212 7636 192484 7664
rect 50212 7624 50218 7636
rect 192478 7624 192484 7636
rect 192536 7624 192542 7676
rect 192570 7624 192576 7676
rect 192628 7664 192634 7676
rect 232038 7664 232044 7676
rect 192628 7636 232044 7664
rect 192628 7624 192634 7636
rect 232038 7624 232044 7636
rect 232096 7624 232102 7676
rect 269942 7624 269948 7676
rect 270000 7664 270006 7676
rect 416682 7664 416688 7676
rect 270000 7636 416688 7664
rect 270000 7624 270006 7636
rect 416682 7624 416688 7636
rect 416740 7624 416746 7676
rect 26510 7556 26516 7608
rect 26568 7596 26574 7608
rect 204346 7596 204352 7608
rect 26568 7568 204352 7596
rect 26568 7556 26574 7568
rect 204346 7556 204352 7568
rect 204404 7556 204410 7608
rect 209774 7556 209780 7608
rect 209832 7596 209838 7608
rect 235074 7596 235080 7608
rect 209832 7568 235080 7596
rect 209832 7556 209838 7568
rect 235074 7556 235080 7568
rect 235132 7556 235138 7608
rect 249978 7556 249984 7608
rect 250036 7596 250042 7608
rect 258442 7596 258448 7608
rect 250036 7568 258448 7596
rect 250036 7556 250042 7568
rect 258442 7556 258448 7568
rect 258500 7556 258506 7608
rect 274082 7556 274088 7608
rect 274140 7596 274146 7608
rect 441522 7596 441528 7608
rect 274140 7568 441528 7596
rect 274140 7556 274146 7568
rect 441522 7556 441528 7568
rect 441580 7556 441586 7608
rect 448606 7556 448612 7608
rect 448664 7596 448670 7608
rect 449802 7596 449808 7608
rect 448664 7568 449808 7596
rect 448664 7556 448670 7568
rect 449802 7556 449808 7568
rect 449860 7556 449866 7608
rect 135254 7488 135260 7540
rect 135312 7528 135318 7540
rect 146938 7528 146944 7540
rect 135312 7500 146944 7528
rect 135312 7488 135318 7500
rect 146938 7488 146944 7500
rect 146996 7488 147002 7540
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 26878 6848 26884 6860
rect 3476 6820 26884 6848
rect 3476 6808 3482 6820
rect 26878 6808 26884 6820
rect 26936 6808 26942 6860
rect 249334 6672 249340 6724
rect 249392 6712 249398 6724
rect 287790 6712 287796 6724
rect 249392 6684 287796 6712
rect 249392 6672 249398 6684
rect 287790 6672 287796 6684
rect 287848 6672 287854 6724
rect 194410 6604 194416 6656
rect 194468 6644 194474 6656
rect 232222 6644 232228 6656
rect 194468 6616 232228 6644
rect 194468 6604 194474 6616
rect 232222 6604 232228 6616
rect 232280 6604 232286 6656
rect 255130 6604 255136 6656
rect 255188 6644 255194 6656
rect 324406 6644 324412 6656
rect 255188 6616 324412 6644
rect 255188 6604 255194 6616
rect 324406 6604 324412 6616
rect 324464 6604 324470 6656
rect 190822 6536 190828 6588
rect 190880 6576 190886 6588
rect 232406 6576 232412 6588
rect 190880 6548 232412 6576
rect 190880 6536 190886 6548
rect 232406 6536 232412 6548
rect 232464 6536 232470 6588
rect 254762 6536 254768 6588
rect 254820 6576 254826 6588
rect 327994 6576 328000 6588
rect 254820 6548 328000 6576
rect 254820 6536 254826 6548
rect 327994 6536 328000 6548
rect 328052 6536 328058 6588
rect 352834 6576 352840 6588
rect 349724 6548 352840 6576
rect 134150 6468 134156 6520
rect 134208 6508 134214 6520
rect 134208 6480 134656 6508
rect 134208 6468 134214 6480
rect 85666 6400 85672 6452
rect 85724 6440 85730 6452
rect 134518 6440 134524 6452
rect 85724 6412 134524 6440
rect 85724 6400 85730 6412
rect 134518 6400 134524 6412
rect 134576 6400 134582 6452
rect 134628 6440 134656 6480
rect 137646 6468 137652 6520
rect 137704 6508 137710 6520
rect 222286 6508 222292 6520
rect 137704 6480 222292 6508
rect 137704 6468 137710 6480
rect 222286 6468 222292 6480
rect 222344 6468 222350 6520
rect 259178 6468 259184 6520
rect 259236 6508 259242 6520
rect 345750 6508 345756 6520
rect 259236 6480 345756 6508
rect 259236 6468 259242 6480
rect 345750 6468 345756 6480
rect 345808 6468 345814 6520
rect 222654 6440 222660 6452
rect 134628 6412 222660 6440
rect 222654 6400 222660 6412
rect 222712 6400 222718 6452
rect 260282 6400 260288 6452
rect 260340 6440 260346 6452
rect 349724 6440 349752 6548
rect 352834 6536 352840 6548
rect 352892 6536 352898 6588
rect 356330 6508 356336 6520
rect 260340 6412 349752 6440
rect 349816 6480 356336 6508
rect 260340 6400 260346 6412
rect 65610 6332 65616 6384
rect 65668 6372 65674 6384
rect 209958 6372 209964 6384
rect 65668 6344 209964 6372
rect 65668 6332 65674 6344
rect 209958 6332 209964 6344
rect 210016 6332 210022 6384
rect 260558 6332 260564 6384
rect 260616 6372 260622 6384
rect 349816 6372 349844 6480
rect 356330 6468 356336 6480
rect 356388 6468 356394 6520
rect 352558 6400 352564 6452
rect 352616 6440 352622 6452
rect 418982 6440 418988 6452
rect 352616 6412 418988 6440
rect 352616 6400 352622 6412
rect 418982 6400 418988 6412
rect 419040 6400 419046 6452
rect 359918 6372 359924 6384
rect 260616 6344 349844 6372
rect 354646 6344 359924 6372
rect 260616 6332 260622 6344
rect 62022 6264 62028 6316
rect 62080 6304 62086 6316
rect 210694 6304 210700 6316
rect 62080 6276 210700 6304
rect 62080 6264 62086 6276
rect 210694 6264 210700 6276
rect 210752 6264 210758 6316
rect 215662 6264 215668 6316
rect 215720 6304 215726 6316
rect 236270 6304 236276 6316
rect 215720 6276 236276 6304
rect 215720 6264 215726 6276
rect 236270 6264 236276 6276
rect 236328 6264 236334 6316
rect 260374 6264 260380 6316
rect 260432 6304 260438 6316
rect 354646 6304 354674 6344
rect 359918 6332 359924 6344
rect 359976 6332 359982 6384
rect 426158 6372 426164 6384
rect 412606 6344 426164 6372
rect 260432 6276 354674 6304
rect 260432 6264 260438 6276
rect 359458 6264 359464 6316
rect 359516 6304 359522 6316
rect 412606 6304 412634 6344
rect 426158 6332 426164 6344
rect 426216 6332 426222 6384
rect 359516 6276 412634 6304
rect 359516 6264 359522 6276
rect 425698 6264 425704 6316
rect 425756 6304 425762 6316
rect 447410 6304 447416 6316
rect 425756 6276 447416 6304
rect 425756 6264 425762 6276
rect 447410 6264 447416 6276
rect 447468 6264 447474 6316
rect 447778 6264 447784 6316
rect 447836 6304 447842 6316
rect 475746 6304 475752 6316
rect 447836 6276 475752 6304
rect 447836 6264 447842 6276
rect 475746 6264 475752 6276
rect 475804 6264 475810 6316
rect 38378 6196 38384 6248
rect 38436 6236 38442 6248
rect 195238 6236 195244 6248
rect 38436 6208 195244 6236
rect 38436 6196 38442 6208
rect 195238 6196 195244 6208
rect 195296 6196 195302 6248
rect 212166 6196 212172 6248
rect 212224 6236 212230 6248
rect 235626 6236 235632 6248
rect 212224 6208 235632 6236
rect 212224 6196 212230 6208
rect 235626 6196 235632 6208
rect 235684 6196 235690 6248
rect 250714 6196 250720 6248
rect 250772 6236 250778 6248
rect 297266 6236 297272 6248
rect 250772 6208 297272 6236
rect 250772 6196 250778 6208
rect 297266 6196 297272 6208
rect 297324 6196 297330 6248
rect 307018 6196 307024 6248
rect 307076 6236 307082 6248
rect 472250 6236 472256 6248
rect 307076 6208 472256 6236
rect 307076 6196 307082 6208
rect 472250 6196 472256 6208
rect 472308 6196 472314 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 200574 6168 200580 6180
rect 4120 6140 200580 6168
rect 4120 6128 4126 6140
rect 200574 6128 200580 6140
rect 200632 6128 200638 6180
rect 208578 6128 208584 6180
rect 208636 6168 208642 6180
rect 234982 6168 234988 6180
rect 208636 6140 234988 6168
rect 208636 6128 208642 6140
rect 234982 6128 234988 6140
rect 235040 6128 235046 6180
rect 249242 6128 249248 6180
rect 249300 6168 249306 6180
rect 291378 6168 291384 6180
rect 249300 6140 291384 6168
rect 249300 6128 249306 6140
rect 291378 6128 291384 6140
rect 291436 6128 291442 6180
rect 292114 6128 292120 6180
rect 292172 6168 292178 6180
rect 543182 6168 543188 6180
rect 292172 6140 543188 6168
rect 292172 6128 292178 6140
rect 543182 6128 543188 6140
rect 543240 6128 543246 6180
rect 234614 5516 234620 5568
rect 234672 5556 234678 5568
rect 239030 5556 239036 5568
rect 234672 5528 239036 5556
rect 234672 5516 234678 5528
rect 239030 5516 239036 5528
rect 239088 5516 239094 5568
rect 124858 5284 124864 5296
rect 103486 5256 124864 5284
rect 24210 5176 24216 5228
rect 24268 5216 24274 5228
rect 98638 5216 98644 5228
rect 24268 5188 98644 5216
rect 24268 5176 24274 5188
rect 98638 5176 98644 5188
rect 98696 5176 98702 5228
rect 99834 5176 99840 5228
rect 99892 5216 99898 5228
rect 103486 5216 103514 5256
rect 124858 5244 124864 5256
rect 124916 5244 124922 5296
rect 99892 5188 103514 5216
rect 99892 5176 99898 5188
rect 245378 5176 245384 5228
rect 245436 5216 245442 5228
rect 265342 5216 265348 5228
rect 245436 5188 265348 5216
rect 245436 5176 245442 5188
rect 265342 5176 265348 5188
rect 265400 5176 265406 5228
rect 370498 5176 370504 5228
rect 370556 5216 370562 5228
rect 433242 5216 433248 5228
rect 370556 5188 433248 5216
rect 370556 5176 370562 5188
rect 433242 5176 433248 5188
rect 433300 5176 433306 5228
rect 35986 5108 35992 5160
rect 36044 5148 36050 5160
rect 58618 5148 58624 5160
rect 36044 5120 58624 5148
rect 36044 5108 36050 5120
rect 58618 5108 58624 5120
rect 58676 5108 58682 5160
rect 58710 5108 58716 5160
rect 58768 5148 58774 5160
rect 209866 5148 209872 5160
rect 58768 5120 209872 5148
rect 58768 5108 58774 5120
rect 209866 5108 209872 5120
rect 209924 5108 209930 5160
rect 249150 5108 249156 5160
rect 249208 5148 249214 5160
rect 290182 5148 290188 5160
rect 249208 5120 290188 5148
rect 249208 5108 249214 5120
rect 290182 5108 290188 5120
rect 290240 5108 290246 5160
rect 363598 5108 363604 5160
rect 363656 5148 363662 5160
rect 429654 5148 429660 5160
rect 363656 5120 429660 5148
rect 363656 5108 363662 5120
rect 429654 5108 429660 5120
rect 429712 5108 429718 5160
rect 54938 5040 54944 5092
rect 54996 5080 55002 5092
rect 208946 5080 208952 5092
rect 54996 5052 208952 5080
rect 54996 5040 55002 5052
rect 208946 5040 208952 5052
rect 209004 5040 209010 5092
rect 221550 5040 221556 5092
rect 221608 5080 221614 5092
rect 236454 5080 236460 5092
rect 221608 5052 236460 5080
rect 221608 5040 221614 5052
rect 236454 5040 236460 5052
rect 236512 5040 236518 5092
rect 249610 5040 249616 5092
rect 249668 5080 249674 5092
rect 293678 5080 293684 5092
rect 249668 5052 293684 5080
rect 249668 5040 249674 5052
rect 293678 5040 293684 5052
rect 293736 5040 293742 5092
rect 302878 5040 302884 5092
rect 302936 5080 302942 5092
rect 372890 5080 372896 5092
rect 302936 5052 372896 5080
rect 302936 5040 302942 5052
rect 372890 5040 372896 5052
rect 372948 5040 372954 5092
rect 429838 5040 429844 5092
rect 429896 5080 429902 5092
rect 454494 5080 454500 5092
rect 429896 5052 454500 5080
rect 429896 5040 429902 5052
rect 454494 5040 454500 5052
rect 454552 5040 454558 5092
rect 47854 4972 47860 5024
rect 47912 5012 47918 5024
rect 207290 5012 207296 5024
rect 47912 4984 207296 5012
rect 47912 4972 47918 4984
rect 207290 4972 207296 4984
rect 207348 4972 207354 5024
rect 218054 4972 218060 5024
rect 218112 5012 218118 5024
rect 236638 5012 236644 5024
rect 218112 4984 236644 5012
rect 218112 4972 218118 4984
rect 236638 4972 236644 4984
rect 236696 4972 236702 5024
rect 245286 4972 245292 5024
rect 245344 5012 245350 5024
rect 268838 5012 268844 5024
rect 245344 4984 268844 5012
rect 245344 4972 245350 4984
rect 268838 4972 268844 4984
rect 268896 4972 268902 5024
rect 271230 4972 271236 5024
rect 271288 5012 271294 5024
rect 415486 5012 415492 5024
rect 271288 4984 415492 5012
rect 271288 4972 271294 4984
rect 415486 4972 415492 4984
rect 415544 4972 415550 5024
rect 450538 4972 450544 5024
rect 450596 5012 450602 5024
rect 582190 5012 582196 5024
rect 450596 4984 582196 5012
rect 450596 4972 450602 4984
rect 582190 4972 582196 4984
rect 582248 4972 582254 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 200390 4944 200396 4956
rect 2924 4916 200396 4944
rect 2924 4904 2930 4916
rect 200390 4904 200396 4916
rect 200448 4904 200454 4956
rect 214466 4904 214472 4956
rect 214524 4944 214530 4956
rect 236178 4944 236184 4956
rect 214524 4916 236184 4944
rect 214524 4904 214530 4916
rect 236178 4904 236184 4916
rect 236236 4904 236242 4956
rect 246482 4904 246488 4956
rect 246540 4944 246546 4956
rect 276014 4944 276020 4956
rect 246540 4916 276020 4944
rect 246540 4904 246546 4916
rect 276014 4904 276020 4916
rect 276072 4904 276078 4956
rect 285214 4904 285220 4956
rect 285272 4944 285278 4956
rect 504174 4944 504180 4956
rect 285272 4916 504180 4944
rect 285272 4904 285278 4916
rect 504174 4904 504180 4916
rect 504232 4904 504238 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 200298 4876 200304 4888
rect 1728 4848 200304 4876
rect 1728 4836 1734 4848
rect 200298 4836 200304 4848
rect 200356 4836 200362 4888
rect 210970 4836 210976 4888
rect 211028 4876 211034 4888
rect 235534 4876 235540 4888
rect 211028 4848 235540 4876
rect 211028 4836 211034 4848
rect 235534 4836 235540 4848
rect 235592 4836 235598 4888
rect 249518 4836 249524 4888
rect 249576 4876 249582 4888
rect 288986 4876 288992 4888
rect 249576 4848 288992 4876
rect 249576 4836 249582 4848
rect 288986 4836 288992 4848
rect 289044 4836 289050 4888
rect 289354 4836 289360 4888
rect 289412 4876 289418 4888
rect 529014 4876 529020 4888
rect 289412 4848 529020 4876
rect 289412 4836 289418 4848
rect 529014 4836 529020 4848
rect 529072 4836 529078 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 200114 4808 200120 4820
rect 624 4780 200120 4808
rect 624 4768 630 4780
rect 200114 4768 200120 4780
rect 200172 4768 200178 4820
rect 207382 4768 207388 4820
rect 207440 4808 207446 4820
rect 234798 4808 234804 4820
rect 207440 4780 234804 4808
rect 207440 4768 207446 4780
rect 234798 4768 234804 4780
rect 234856 4768 234862 4820
rect 249426 4768 249432 4820
rect 249484 4808 249490 4820
rect 292574 4808 292580 4820
rect 249484 4780 292580 4808
rect 249484 4768 249490 4780
rect 292574 4768 292580 4780
rect 292632 4768 292638 4820
rect 294782 4768 294788 4820
rect 294840 4808 294846 4820
rect 558546 4808 558552 4820
rect 294840 4780 558552 4808
rect 294840 4768 294846 4780
rect 558546 4768 558552 4780
rect 558604 4768 558610 4820
rect 84028 4168 84194 4196
rect 60826 4088 60832 4140
rect 60884 4128 60890 4140
rect 71038 4128 71044 4140
rect 60884 4100 71044 4128
rect 60884 4088 60890 4100
rect 71038 4088 71044 4100
rect 71096 4088 71102 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 80698 4128 80704 4140
rect 73856 4100 80704 4128
rect 73856 4088 73862 4100
rect 80698 4088 80704 4100
rect 80756 4088 80762 4140
rect 82078 4088 82084 4140
rect 82136 4128 82142 4140
rect 84028 4128 84056 4168
rect 82136 4100 84056 4128
rect 84166 4128 84194 4168
rect 124674 4156 124680 4208
rect 124732 4196 124738 4208
rect 126238 4196 126244 4208
rect 124732 4168 126244 4196
rect 124732 4156 124738 4168
rect 126238 4156 126244 4168
rect 126296 4156 126302 4208
rect 241238 4156 241244 4208
rect 241296 4196 241302 4208
rect 242894 4196 242900 4208
rect 241296 4168 242900 4196
rect 241296 4156 241302 4168
rect 242894 4156 242900 4168
rect 242952 4156 242958 4208
rect 93118 4128 93124 4140
rect 84166 4100 93124 4128
rect 82136 4088 82142 4100
rect 93118 4088 93124 4100
rect 93176 4088 93182 4140
rect 146938 4088 146944 4140
rect 146996 4128 147002 4140
rect 223574 4128 223580 4140
rect 146996 4100 223580 4128
rect 146996 4088 147002 4100
rect 223574 4088 223580 4100
rect 223632 4088 223638 4140
rect 228726 4088 228732 4140
rect 228784 4128 228790 4140
rect 237650 4128 237656 4140
rect 228784 4100 237656 4128
rect 228784 4088 228790 4100
rect 237650 4088 237656 4100
rect 237708 4088 237714 4140
rect 257338 4088 257344 4140
rect 257396 4128 257402 4140
rect 258258 4128 258264 4140
rect 257396 4100 258264 4128
rect 257396 4088 257402 4100
rect 258258 4088 258264 4100
rect 258316 4088 258322 4140
rect 353938 4088 353944 4140
rect 353996 4128 354002 4140
rect 355226 4128 355232 4140
rect 353996 4100 355232 4128
rect 353996 4088 354002 4100
rect 355226 4088 355232 4100
rect 355284 4088 355290 4140
rect 410518 4088 410524 4140
rect 410576 4128 410582 4140
rect 424962 4128 424968 4140
rect 410576 4100 424968 4128
rect 410576 4088 410582 4100
rect 424962 4088 424968 4100
rect 425020 4088 425026 4140
rect 453298 4088 453304 4140
rect 453356 4128 453362 4140
rect 455690 4128 455696 4140
rect 453356 4100 455696 4128
rect 453356 4088 453362 4100
rect 455690 4088 455696 4100
rect 455748 4088 455754 4140
rect 460198 4088 460204 4140
rect 460256 4128 460262 4140
rect 462774 4128 462780 4140
rect 460256 4100 462780 4128
rect 460256 4088 460262 4100
rect 462774 4088 462780 4100
rect 462832 4088 462838 4140
rect 479518 4088 479524 4140
rect 479576 4128 479582 4140
rect 480530 4128 480536 4140
rect 479576 4100 480536 4128
rect 479576 4088 479582 4100
rect 480530 4088 480536 4100
rect 480588 4088 480594 4140
rect 518158 4088 518164 4140
rect 518216 4128 518222 4140
rect 520734 4128 520740 4140
rect 518216 4100 520740 4128
rect 518216 4088 518222 4100
rect 520734 4088 520740 4100
rect 520792 4088 520798 4140
rect 565078 4088 565084 4140
rect 565136 4128 565142 4140
rect 568022 4128 568028 4140
rect 565136 4100 568028 4128
rect 565136 4088 565142 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 46198 4060 46204 4072
rect 34848 4032 46204 4060
rect 34848 4020 34854 4032
rect 46198 4020 46204 4032
rect 46256 4020 46262 4072
rect 57238 4020 57244 4072
rect 57296 4060 57302 4072
rect 87598 4060 87604 4072
rect 57296 4032 87604 4060
rect 57296 4020 57302 4032
rect 87598 4020 87604 4032
rect 87656 4020 87662 4072
rect 101030 4020 101036 4072
rect 101088 4060 101094 4072
rect 104158 4060 104164 4072
rect 101088 4032 104164 4060
rect 101088 4020 101094 4032
rect 104158 4020 104164 4032
rect 104216 4020 104222 4072
rect 122098 4060 122104 4072
rect 113146 4032 122104 4060
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 35158 3992 35164 4004
rect 19484 3964 35164 3992
rect 19484 3952 19490 3964
rect 35158 3952 35164 3964
rect 35216 3952 35222 4004
rect 56042 3952 56048 4004
rect 56100 3992 56106 4004
rect 65518 3992 65524 4004
rect 56100 3964 65524 3992
rect 56100 3952 56106 3964
rect 65518 3952 65524 3964
rect 65576 3952 65582 4004
rect 71498 3952 71504 4004
rect 71556 3992 71562 4004
rect 101398 3992 101404 4004
rect 71556 3964 101404 3992
rect 71556 3952 71562 3964
rect 101398 3952 101404 3964
rect 101456 3952 101462 4004
rect 103330 3952 103336 4004
rect 103388 3992 103394 4004
rect 113146 3992 113174 4032
rect 122098 4020 122104 4032
rect 122156 4020 122162 4072
rect 129366 4020 129372 4072
rect 129424 4060 129430 4072
rect 221090 4060 221096 4072
rect 129424 4032 221096 4060
rect 129424 4020 129430 4032
rect 221090 4020 221096 4032
rect 221148 4020 221154 4072
rect 238202 4060 238208 4072
rect 229664 4032 238208 4060
rect 103388 3964 113174 3992
rect 103388 3952 103394 3964
rect 117590 3952 117596 4004
rect 117648 3992 117654 4004
rect 214558 3992 214564 4004
rect 117648 3964 214564 3992
rect 117648 3952 117654 3964
rect 214558 3952 214564 3964
rect 214616 3952 214622 4004
rect 223758 3952 223764 4004
rect 223816 3992 223822 4004
rect 228358 3992 228364 4004
rect 223816 3964 228364 3992
rect 223816 3952 223822 3964
rect 228358 3952 228364 3964
rect 228416 3952 228422 4004
rect 28902 3884 28908 3936
rect 28960 3924 28966 3936
rect 47578 3924 47584 3936
rect 28960 3896 47584 3924
rect 28960 3884 28966 3896
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 53742 3884 53748 3936
rect 53800 3924 53806 3936
rect 88978 3924 88984 3936
rect 53800 3896 88984 3924
rect 53800 3884 53806 3896
rect 88978 3884 88984 3896
rect 89036 3884 89042 3936
rect 92750 3884 92756 3936
rect 92808 3924 92814 3936
rect 97258 3924 97264 3936
rect 92808 3896 97264 3924
rect 92808 3884 92814 3896
rect 97258 3884 97264 3896
rect 97316 3884 97322 3936
rect 112806 3884 112812 3936
rect 112864 3924 112870 3936
rect 116578 3924 116584 3936
rect 112864 3896 116584 3924
rect 112864 3884 112870 3896
rect 116578 3884 116584 3896
rect 116636 3884 116642 3936
rect 121086 3884 121092 3936
rect 121144 3924 121150 3936
rect 220078 3924 220084 3936
rect 121144 3896 220084 3924
rect 121144 3884 121150 3896
rect 220078 3884 220084 3896
rect 220136 3884 220142 3936
rect 226334 3884 226340 3936
rect 226392 3924 226398 3936
rect 229664 3924 229692 4032
rect 238202 4020 238208 4032
rect 238260 4020 238266 4072
rect 256142 4020 256148 4072
rect 256200 4060 256206 4072
rect 260650 4060 260656 4072
rect 256200 4032 260656 4060
rect 256200 4020 256206 4032
rect 260650 4020 260656 4032
rect 260708 4020 260714 4072
rect 406378 4020 406384 4072
rect 406436 4060 406442 4072
rect 406436 4032 412634 4060
rect 406436 4020 406442 4032
rect 259270 3952 259276 4004
rect 259328 3992 259334 4004
rect 266722 3992 266728 4004
rect 259328 3964 266728 3992
rect 259328 3952 259334 3964
rect 266722 3952 266728 3964
rect 266780 3952 266786 4004
rect 266998 3952 267004 4004
rect 267056 3992 267062 4004
rect 271230 3992 271236 4004
rect 267056 3964 271236 3992
rect 267056 3952 267062 3964
rect 271230 3952 271236 3964
rect 271288 3952 271294 4004
rect 273898 3952 273904 4004
rect 273956 3992 273962 4004
rect 278314 3992 278320 4004
rect 273956 3964 278320 3992
rect 273956 3952 273962 3964
rect 278314 3952 278320 3964
rect 278372 3952 278378 4004
rect 296070 3952 296076 4004
rect 296128 3992 296134 4004
rect 298186 3992 298192 4004
rect 296128 3964 298192 3992
rect 296128 3952 296134 3964
rect 298186 3952 298192 3964
rect 298244 3952 298250 4004
rect 392670 3952 392676 4004
rect 392728 3992 392734 4004
rect 394234 3992 394240 4004
rect 392728 3964 394240 3992
rect 392728 3952 392734 3964
rect 394234 3952 394240 3964
rect 394292 3952 394298 4004
rect 412606 3992 412634 4032
rect 418798 4020 418804 4072
rect 418856 4060 418862 4072
rect 436738 4060 436744 4072
rect 418856 4032 436744 4060
rect 418856 4020 418862 4032
rect 436738 4020 436744 4032
rect 436796 4020 436802 4072
rect 464338 4020 464344 4072
rect 464396 4060 464402 4072
rect 473446 4060 473452 4072
rect 464396 4032 473452 4060
rect 464396 4020 464402 4032
rect 473446 4020 473452 4032
rect 473504 4020 473510 4072
rect 432046 3992 432052 4004
rect 412606 3964 432052 3992
rect 432046 3952 432052 3964
rect 432104 3952 432110 4004
rect 436830 3952 436836 4004
rect 436888 3992 436894 4004
rect 436888 3964 447134 3992
rect 436888 3952 436894 3964
rect 237926 3924 237932 3936
rect 226392 3896 229692 3924
rect 229848 3896 237932 3924
rect 226392 3884 226398 3896
rect 11146 3816 11152 3868
rect 11204 3856 11210 3868
rect 28258 3856 28264 3868
rect 11204 3828 28264 3856
rect 11204 3816 11210 3828
rect 28258 3816 28264 3828
rect 28316 3816 28322 3868
rect 46658 3816 46664 3868
rect 46716 3856 46722 3868
rect 94498 3856 94504 3868
rect 46716 3828 94504 3856
rect 46716 3816 46722 3828
rect 94498 3816 94504 3828
rect 94556 3816 94562 3868
rect 96246 3816 96252 3868
rect 96304 3856 96310 3868
rect 210418 3856 210424 3868
rect 96304 3828 210424 3856
rect 96304 3816 96310 3828
rect 210418 3816 210424 3828
rect 210476 3816 210482 3868
rect 225138 3816 225144 3868
rect 225196 3856 225202 3868
rect 229848 3856 229876 3896
rect 237926 3884 237932 3896
rect 237984 3884 237990 3936
rect 256050 3884 256056 3936
rect 256108 3924 256114 3936
rect 267734 3924 267740 3936
rect 256108 3896 267740 3924
rect 256108 3884 256114 3896
rect 267734 3884 267740 3896
rect 267792 3884 267798 3936
rect 304258 3884 304264 3936
rect 304316 3924 304322 3936
rect 351638 3924 351644 3936
rect 304316 3896 351644 3924
rect 304316 3884 304322 3896
rect 351638 3884 351644 3896
rect 351696 3884 351702 3936
rect 407758 3884 407764 3936
rect 407816 3924 407822 3936
rect 435542 3924 435548 3936
rect 407816 3896 435548 3924
rect 407816 3884 407822 3896
rect 435542 3884 435548 3896
rect 435600 3884 435606 3936
rect 225196 3828 229876 3856
rect 225196 3816 225202 3828
rect 229922 3816 229928 3868
rect 229980 3856 229986 3868
rect 238110 3856 238116 3868
rect 229980 3828 238116 3856
rect 229980 3816 229986 3828
rect 238110 3816 238116 3828
rect 238168 3816 238174 3868
rect 242802 3816 242808 3868
rect 242860 3856 242866 3868
rect 251174 3856 251180 3868
rect 242860 3828 251180 3856
rect 242860 3816 242866 3828
rect 251174 3816 251180 3828
rect 251232 3816 251238 3868
rect 255958 3816 255964 3868
rect 256016 3856 256022 3868
rect 259454 3856 259460 3868
rect 256016 3828 259460 3856
rect 256016 3816 256022 3828
rect 259454 3816 259460 3828
rect 259512 3816 259518 3868
rect 261478 3816 261484 3868
rect 261536 3856 261542 3868
rect 277118 3856 277124 3868
rect 261536 3828 277124 3856
rect 261536 3816 261542 3828
rect 277118 3816 277124 3828
rect 277176 3816 277182 3868
rect 299566 3816 299572 3868
rect 299624 3856 299630 3868
rect 300762 3856 300768 3868
rect 299624 3828 300768 3856
rect 299624 3816 299630 3828
rect 300762 3816 300768 3828
rect 300820 3816 300826 3868
rect 322198 3816 322204 3868
rect 322256 3856 322262 3868
rect 383562 3856 383568 3868
rect 322256 3828 383568 3856
rect 322256 3816 322262 3828
rect 383562 3816 383568 3828
rect 383620 3816 383626 3868
rect 393958 3816 393964 3868
rect 394016 3856 394022 3868
rect 422570 3856 422576 3868
rect 394016 3828 422576 3856
rect 394016 3816 394022 3828
rect 422570 3816 422576 3828
rect 422628 3816 422634 3868
rect 440878 3816 440884 3868
rect 440936 3856 440942 3868
rect 445018 3856 445024 3868
rect 440936 3828 445024 3856
rect 440936 3816 440942 3828
rect 445018 3816 445024 3828
rect 445076 3816 445082 3868
rect 447106 3856 447134 3964
rect 476758 3952 476764 4004
rect 476816 3992 476822 4004
rect 485222 3992 485228 4004
rect 476816 3964 485228 3992
rect 476816 3952 476822 3964
rect 485222 3952 485228 3964
rect 485280 3952 485286 4004
rect 472618 3884 472624 3936
rect 472676 3924 472682 3936
rect 491110 3924 491116 3936
rect 472676 3896 491116 3924
rect 472676 3884 472682 3896
rect 491110 3884 491116 3896
rect 491168 3884 491174 3936
rect 461578 3856 461584 3868
rect 447106 3828 461584 3856
rect 461578 3816 461584 3828
rect 461636 3816 461642 3868
rect 468478 3816 468484 3868
rect 468536 3856 468542 3868
rect 498194 3856 498200 3868
rect 468536 3828 498200 3856
rect 468536 3816 468542 3828
rect 498194 3816 498200 3828
rect 498252 3816 498258 3868
rect 503070 3816 503076 3868
rect 503128 3856 503134 3868
rect 530118 3856 530124 3868
rect 503128 3828 530124 3856
rect 503128 3816 503134 3828
rect 530118 3816 530124 3828
rect 530176 3816 530182 3868
rect 20622 3748 20628 3800
rect 20680 3788 20686 3800
rect 39298 3788 39304 3800
rect 20680 3760 39304 3788
rect 20680 3748 20686 3760
rect 39298 3748 39304 3760
rect 39356 3748 39362 3800
rect 45370 3748 45376 3800
rect 45428 3788 45434 3800
rect 57146 3788 57152 3800
rect 45428 3760 57152 3788
rect 45428 3748 45434 3760
rect 57146 3748 57152 3760
rect 57204 3748 57210 3800
rect 63218 3748 63224 3800
rect 63276 3788 63282 3800
rect 210142 3788 210148 3800
rect 63276 3760 210148 3788
rect 63276 3748 63282 3760
rect 210142 3748 210148 3760
rect 210200 3748 210206 3800
rect 219250 3748 219256 3800
rect 219308 3788 219314 3800
rect 231118 3788 231124 3800
rect 219308 3760 231124 3788
rect 219308 3748 219314 3760
rect 231118 3748 231124 3760
rect 231176 3748 231182 3800
rect 252002 3748 252008 3800
rect 252060 3788 252066 3800
rect 252060 3760 258074 3788
rect 252060 3748 252066 3760
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 36538 3720 36544 3732
rect 13596 3692 36544 3720
rect 13596 3680 13602 3692
rect 36538 3680 36544 3692
rect 36596 3680 36602 3732
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 50338 3720 50344 3732
rect 41932 3692 50344 3720
rect 41932 3680 41938 3692
rect 50338 3680 50344 3692
rect 50396 3680 50402 3732
rect 51350 3680 51356 3732
rect 51408 3720 51414 3732
rect 208762 3720 208768 3732
rect 51408 3692 208768 3720
rect 51408 3680 51414 3692
rect 208762 3680 208768 3692
rect 208820 3680 208826 3732
rect 216858 3680 216864 3732
rect 216916 3720 216922 3732
rect 229830 3720 229836 3732
rect 216916 3692 229836 3720
rect 216916 3680 216922 3692
rect 229830 3680 229836 3692
rect 229888 3680 229894 3732
rect 242618 3680 242624 3732
rect 242676 3720 242682 3732
rect 252370 3720 252376 3732
rect 242676 3692 252376 3720
rect 242676 3680 242682 3692
rect 252370 3680 252376 3692
rect 252428 3680 252434 3732
rect 258046 3720 258074 3760
rect 259362 3748 259368 3800
rect 259420 3788 259426 3800
rect 349246 3788 349252 3800
rect 259420 3760 349252 3788
rect 259420 3748 259426 3760
rect 349246 3748 349252 3760
rect 349304 3748 349310 3800
rect 381538 3748 381544 3800
rect 381596 3788 381602 3800
rect 411898 3788 411904 3800
rect 381596 3760 411904 3788
rect 381596 3748 381602 3760
rect 411898 3748 411904 3760
rect 411956 3748 411962 3800
rect 411990 3748 411996 3800
rect 412048 3788 412054 3800
rect 440326 3788 440332 3800
rect 412048 3760 440332 3788
rect 412048 3748 412054 3760
rect 440326 3748 440332 3760
rect 440384 3748 440390 3800
rect 443638 3748 443644 3800
rect 443696 3788 443702 3800
rect 443696 3760 447134 3788
rect 443696 3748 443702 3760
rect 305546 3720 305552 3732
rect 258046 3692 305552 3720
rect 305546 3680 305552 3692
rect 305604 3680 305610 3732
rect 327718 3680 327724 3732
rect 327776 3720 327782 3732
rect 390646 3720 390652 3732
rect 327776 3692 390652 3720
rect 327776 3680 327782 3692
rect 390646 3680 390652 3692
rect 390704 3680 390710 3732
rect 396718 3680 396724 3732
rect 396776 3720 396782 3732
rect 443822 3720 443828 3732
rect 396776 3692 443828 3720
rect 396776 3680 396782 3692
rect 443822 3680 443828 3692
rect 443880 3680 443886 3732
rect 447106 3720 447134 3760
rect 461670 3748 461676 3800
rect 461728 3788 461734 3800
rect 505370 3788 505376 3800
rect 461728 3760 505376 3788
rect 461728 3748 461734 3760
rect 505370 3748 505376 3760
rect 505428 3748 505434 3800
rect 468662 3720 468668 3732
rect 447106 3692 468668 3720
rect 468662 3680 468668 3692
rect 468720 3680 468726 3732
rect 475378 3680 475384 3732
rect 475436 3720 475442 3732
rect 487614 3720 487620 3732
rect 475436 3692 487620 3720
rect 475436 3680 475442 3692
rect 487614 3680 487620 3692
rect 487672 3680 487678 3732
rect 489178 3680 489184 3732
rect 489236 3720 489242 3732
rect 540790 3720 540796 3732
rect 489236 3692 540796 3720
rect 489236 3680 489242 3692
rect 540790 3680 540796 3692
rect 540848 3680 540854 3732
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 21358 3652 21364 3664
rect 10008 3624 21364 3652
rect 10008 3612 10014 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 25314 3612 25320 3664
rect 25372 3652 25378 3664
rect 204254 3652 204260 3664
rect 25372 3624 204260 3652
rect 25372 3612 25378 3624
rect 204254 3612 204260 3624
rect 204312 3612 204318 3664
rect 213362 3612 213368 3664
rect 213420 3652 213426 3664
rect 231210 3652 231216 3664
rect 213420 3624 231216 3652
rect 213420 3612 213426 3624
rect 231210 3612 231216 3624
rect 231268 3612 231274 3664
rect 238110 3612 238116 3664
rect 238168 3652 238174 3664
rect 240962 3652 240968 3664
rect 238168 3624 240968 3652
rect 238168 3612 238174 3624
rect 240962 3612 240968 3624
rect 241020 3612 241026 3664
rect 246298 3612 246304 3664
rect 246356 3652 246362 3664
rect 255866 3652 255872 3664
rect 246356 3624 255872 3652
rect 246356 3612 246362 3624
rect 255866 3612 255872 3624
rect 255924 3612 255930 3664
rect 262950 3652 262956 3664
rect 258046 3624 262956 3652
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 7708 3556 16574 3584
rect 7708 3544 7714 3556
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15838 3516 15844 3528
rect 14792 3488 15844 3516
rect 14792 3476 14798 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16546 3516 16574 3556
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17862 3584 17868 3596
rect 17092 3556 17868 3584
rect 17092 3544 17098 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 19242 3584 19248 3596
rect 18288 3556 19248 3584
rect 18288 3544 18294 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 25498 3584 25504 3596
rect 21876 3556 25504 3584
rect 21876 3544 21882 3556
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 29638 3584 29644 3596
rect 27764 3556 29644 3584
rect 27764 3544 27770 3556
rect 29638 3544 29644 3556
rect 29696 3544 29702 3596
rect 32398 3544 32404 3596
rect 32456 3584 32462 3596
rect 33042 3584 33048 3596
rect 32456 3556 33048 3584
rect 32456 3544 32462 3556
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 40678 3544 40684 3596
rect 40736 3584 40742 3596
rect 41322 3584 41328 3596
rect 40736 3556 41328 3584
rect 40736 3544 40742 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 44082 3584 44088 3596
rect 43128 3556 44088 3584
rect 43128 3544 43134 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45462 3584 45468 3596
rect 44324 3556 45468 3584
rect 44324 3544 44330 3556
rect 45462 3544 45468 3556
rect 45520 3544 45526 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 54478 3584 54484 3596
rect 52604 3556 54484 3584
rect 52604 3544 52610 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64782 3584 64788 3596
rect 64380 3556 64788 3584
rect 64380 3544 64386 3556
rect 64782 3544 64788 3556
rect 64840 3544 64846 3596
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 68922 3584 68928 3596
rect 67968 3556 68928 3584
rect 67968 3544 67974 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 72602 3544 72608 3596
rect 72660 3584 72666 3596
rect 73062 3584 73068 3596
rect 72660 3556 73068 3584
rect 72660 3544 72666 3556
rect 73062 3544 73068 3556
rect 73120 3544 73126 3596
rect 76190 3544 76196 3596
rect 76248 3584 76254 3596
rect 77202 3584 77208 3596
rect 76248 3556 77208 3584
rect 76248 3544 76254 3556
rect 77202 3544 77208 3556
rect 77260 3544 77266 3596
rect 77386 3544 77392 3596
rect 77444 3584 77450 3596
rect 79318 3584 79324 3596
rect 77444 3556 79324 3584
rect 77444 3544 77450 3556
rect 79318 3544 79324 3556
rect 79376 3544 79382 3596
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 84102 3584 84108 3596
rect 83332 3556 84108 3584
rect 83332 3544 83338 3556
rect 84102 3544 84108 3556
rect 84160 3544 84166 3596
rect 84470 3544 84476 3596
rect 84528 3584 84534 3596
rect 85482 3584 85488 3596
rect 84528 3556 85488 3584
rect 84528 3544 84534 3556
rect 85482 3544 85488 3556
rect 85540 3544 85546 3596
rect 89162 3544 89168 3596
rect 89220 3584 89226 3596
rect 90358 3584 90364 3596
rect 89220 3556 90364 3584
rect 89220 3544 89226 3556
rect 90358 3544 90364 3556
rect 90416 3544 90422 3596
rect 91554 3544 91560 3596
rect 91612 3584 91618 3596
rect 92382 3584 92388 3596
rect 91612 3556 92388 3584
rect 91612 3544 91618 3556
rect 92382 3544 92388 3556
rect 92440 3544 92446 3596
rect 98638 3544 98644 3596
rect 98696 3584 98702 3596
rect 99282 3584 99288 3596
rect 98696 3556 99288 3584
rect 98696 3544 98702 3556
rect 99282 3544 99288 3556
rect 99340 3544 99346 3596
rect 102226 3544 102232 3596
rect 102284 3584 102290 3596
rect 103422 3584 103428 3596
rect 102284 3556 103428 3584
rect 102284 3544 102290 3556
rect 103422 3544 103428 3556
rect 103480 3544 103486 3596
rect 105722 3544 105728 3596
rect 105780 3584 105786 3596
rect 106182 3584 106188 3596
rect 105780 3556 106188 3584
rect 105780 3544 105786 3556
rect 106182 3544 106188 3556
rect 106240 3544 106246 3596
rect 106918 3544 106924 3596
rect 106976 3584 106982 3596
rect 107562 3584 107568 3596
rect 106976 3556 107568 3584
rect 106976 3544 106982 3556
rect 107562 3544 107568 3556
rect 107620 3544 107626 3596
rect 108114 3544 108120 3596
rect 108172 3584 108178 3596
rect 108942 3584 108948 3596
rect 108172 3556 108948 3584
rect 108172 3544 108178 3556
rect 108942 3544 108948 3556
rect 109000 3544 109006 3596
rect 109310 3544 109316 3596
rect 109368 3584 109374 3596
rect 111058 3584 111064 3596
rect 109368 3556 111064 3584
rect 109368 3544 109374 3556
rect 111058 3544 111064 3556
rect 111116 3544 111122 3596
rect 111610 3544 111616 3596
rect 111668 3584 111674 3596
rect 112438 3584 112444 3596
rect 111668 3556 112444 3584
rect 111668 3544 111674 3556
rect 112438 3544 112444 3556
rect 112496 3544 112502 3596
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 115198 3584 115204 3596
rect 114060 3556 115204 3584
rect 114060 3544 114066 3556
rect 115198 3544 115204 3556
rect 115256 3544 115262 3596
rect 116394 3544 116400 3596
rect 116452 3584 116458 3596
rect 117222 3584 117228 3596
rect 116452 3556 117228 3584
rect 116452 3544 116458 3556
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 124122 3584 124128 3596
rect 123536 3556 124128 3584
rect 123536 3544 123542 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 125870 3544 125876 3596
rect 125928 3584 125934 3596
rect 126882 3584 126888 3596
rect 125928 3556 126888 3584
rect 125928 3544 125934 3556
rect 126882 3544 126888 3556
rect 126940 3544 126946 3596
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 128262 3584 128268 3596
rect 127032 3556 128268 3584
rect 127032 3544 127038 3556
rect 128262 3544 128268 3556
rect 128320 3544 128326 3596
rect 130562 3544 130568 3596
rect 130620 3584 130626 3596
rect 131022 3584 131028 3596
rect 130620 3556 131028 3584
rect 130620 3544 130626 3556
rect 131022 3544 131028 3556
rect 131080 3544 131086 3596
rect 132954 3544 132960 3596
rect 133012 3584 133018 3596
rect 133782 3584 133788 3596
rect 133012 3556 133788 3584
rect 133012 3544 133018 3556
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 136450 3544 136456 3596
rect 136508 3584 136514 3596
rect 137278 3584 137284 3596
rect 136508 3556 137284 3584
rect 136508 3544 136514 3556
rect 137278 3544 137284 3556
rect 137336 3544 137342 3596
rect 140038 3544 140044 3596
rect 140096 3584 140102 3596
rect 146938 3584 146944 3596
rect 140096 3556 146944 3584
rect 140096 3544 140102 3556
rect 146938 3544 146944 3556
rect 146996 3544 147002 3596
rect 147122 3544 147128 3596
rect 147180 3584 147186 3596
rect 147582 3584 147588 3596
rect 147180 3556 147588 3584
rect 147180 3544 147186 3556
rect 147582 3544 147588 3556
rect 147640 3544 147646 3596
rect 148318 3544 148324 3596
rect 148376 3584 148382 3596
rect 148962 3584 148968 3596
rect 148376 3556 148968 3584
rect 148376 3544 148382 3556
rect 148962 3544 148968 3556
rect 149020 3544 149026 3596
rect 149514 3544 149520 3596
rect 149572 3584 149578 3596
rect 150342 3584 150348 3596
rect 149572 3556 150348 3584
rect 149572 3544 149578 3556
rect 150342 3544 150348 3556
rect 150400 3544 150406 3596
rect 151814 3544 151820 3596
rect 151872 3584 151878 3596
rect 153102 3584 153108 3596
rect 151872 3556 153108 3584
rect 151872 3544 151878 3556
rect 153102 3544 153108 3556
rect 153160 3544 153166 3596
rect 154206 3544 154212 3596
rect 154264 3584 154270 3596
rect 155218 3584 155224 3596
rect 154264 3556 155224 3584
rect 154264 3544 154270 3556
rect 155218 3544 155224 3556
rect 155276 3544 155282 3596
rect 155402 3544 155408 3596
rect 155460 3584 155466 3596
rect 155862 3584 155868 3596
rect 155460 3556 155868 3584
rect 155460 3544 155466 3556
rect 155862 3544 155868 3556
rect 155920 3544 155926 3596
rect 156598 3544 156604 3596
rect 156656 3584 156662 3596
rect 157242 3584 157248 3596
rect 156656 3556 157248 3584
rect 156656 3544 156662 3556
rect 157242 3544 157248 3556
rect 157300 3544 157306 3596
rect 157794 3544 157800 3596
rect 157852 3584 157858 3596
rect 158622 3584 158628 3596
rect 157852 3556 158628 3584
rect 157852 3544 157858 3556
rect 158622 3544 158628 3556
rect 158680 3544 158686 3596
rect 158898 3544 158904 3596
rect 158956 3584 158962 3596
rect 160002 3584 160008 3596
rect 158956 3556 160008 3584
rect 158956 3544 158962 3556
rect 160002 3544 160008 3556
rect 160060 3544 160066 3596
rect 160094 3544 160100 3596
rect 160152 3584 160158 3596
rect 161198 3584 161204 3596
rect 160152 3556 161204 3584
rect 160152 3544 160158 3556
rect 161198 3544 161204 3556
rect 161256 3544 161262 3596
rect 163682 3544 163688 3596
rect 163740 3584 163746 3596
rect 164142 3584 164148 3596
rect 163740 3556 164148 3584
rect 163740 3544 163746 3556
rect 164142 3544 164148 3556
rect 164200 3544 164206 3596
rect 164878 3544 164884 3596
rect 164936 3584 164942 3596
rect 165522 3584 165528 3596
rect 164936 3556 165528 3584
rect 164936 3544 164942 3556
rect 165522 3544 165528 3556
rect 165580 3544 165586 3596
rect 166074 3544 166080 3596
rect 166132 3584 166138 3596
rect 166902 3584 166908 3596
rect 166132 3556 166908 3584
rect 166132 3544 166138 3556
rect 166902 3544 166908 3556
rect 166960 3544 166966 3596
rect 167178 3544 167184 3596
rect 167236 3584 167242 3596
rect 169018 3584 169024 3596
rect 167236 3556 169024 3584
rect 167236 3544 167242 3556
rect 169018 3544 169024 3556
rect 169076 3544 169082 3596
rect 171962 3544 171968 3596
rect 172020 3584 172026 3596
rect 173158 3584 173164 3596
rect 172020 3556 173164 3584
rect 172020 3544 172026 3556
rect 173158 3544 173164 3556
rect 173216 3544 173222 3596
rect 174262 3544 174268 3596
rect 174320 3584 174326 3596
rect 175182 3584 175188 3596
rect 174320 3556 175188 3584
rect 174320 3544 174326 3556
rect 175182 3544 175188 3556
rect 175240 3544 175246 3596
rect 175458 3544 175464 3596
rect 175516 3584 175522 3596
rect 176562 3584 176568 3596
rect 175516 3556 176568 3584
rect 175516 3544 175522 3556
rect 176562 3544 176568 3556
rect 176620 3544 176626 3596
rect 176654 3544 176660 3596
rect 176712 3584 176718 3596
rect 177942 3584 177948 3596
rect 176712 3556 177948 3584
rect 176712 3544 176718 3556
rect 177942 3544 177948 3556
rect 178000 3544 178006 3596
rect 180242 3544 180248 3596
rect 180300 3584 180306 3596
rect 180702 3584 180708 3596
rect 180300 3556 180708 3584
rect 180300 3544 180306 3556
rect 180702 3544 180708 3556
rect 180760 3544 180766 3596
rect 181438 3544 181444 3596
rect 181496 3584 181502 3596
rect 182082 3584 182088 3596
rect 181496 3556 182088 3584
rect 181496 3544 181502 3556
rect 182082 3544 182088 3556
rect 182140 3544 182146 3596
rect 182542 3544 182548 3596
rect 182600 3584 182606 3596
rect 183462 3584 183468 3596
rect 182600 3556 183468 3584
rect 182600 3544 182606 3556
rect 183462 3544 183468 3556
rect 183520 3544 183526 3596
rect 183738 3544 183744 3596
rect 183796 3584 183802 3596
rect 184842 3584 184848 3596
rect 183796 3556 184848 3584
rect 183796 3544 183802 3556
rect 184842 3544 184848 3556
rect 184900 3544 184906 3596
rect 186130 3544 186136 3596
rect 186188 3584 186194 3596
rect 186958 3584 186964 3596
rect 186188 3556 186964 3584
rect 186188 3544 186194 3556
rect 186958 3544 186964 3556
rect 187016 3544 187022 3596
rect 187326 3544 187332 3596
rect 187384 3584 187390 3596
rect 188338 3584 188344 3596
rect 187384 3556 188344 3584
rect 187384 3544 187390 3556
rect 188338 3544 188344 3556
rect 188396 3544 188402 3596
rect 188522 3544 188528 3596
rect 188580 3584 188586 3596
rect 188982 3584 188988 3596
rect 188580 3556 188988 3584
rect 188580 3544 188586 3556
rect 188982 3544 188988 3556
rect 189040 3544 189046 3596
rect 189718 3544 189724 3596
rect 189776 3584 189782 3596
rect 191098 3584 191104 3596
rect 189776 3556 191104 3584
rect 189776 3544 189782 3556
rect 191098 3544 191104 3556
rect 191156 3544 191162 3596
rect 192018 3544 192024 3596
rect 192076 3584 192082 3596
rect 192570 3584 192576 3596
rect 192076 3556 192576 3584
rect 192076 3544 192082 3556
rect 192570 3544 192576 3556
rect 192628 3544 192634 3596
rect 193214 3544 193220 3596
rect 193272 3584 193278 3596
rect 194502 3584 194508 3596
rect 193272 3556 194508 3584
rect 193272 3544 193278 3556
rect 194502 3544 194508 3556
rect 194560 3544 194566 3596
rect 196802 3544 196808 3596
rect 196860 3584 196866 3596
rect 197262 3584 197268 3596
rect 196860 3556 197268 3584
rect 196860 3544 196866 3556
rect 197262 3544 197268 3556
rect 197320 3544 197326 3596
rect 197906 3544 197912 3596
rect 197964 3584 197970 3596
rect 198642 3584 198648 3596
rect 197964 3556 198648 3584
rect 197964 3544 197970 3556
rect 198642 3544 198648 3556
rect 198700 3544 198706 3596
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 223758 3584 223764 3596
rect 201552 3556 223764 3584
rect 201552 3544 201558 3556
rect 223758 3544 223764 3556
rect 223816 3544 223822 3596
rect 235442 3584 235448 3596
rect 223868 3556 235448 3584
rect 200942 3516 200948 3528
rect 16546 3488 200948 3516
rect 200942 3476 200948 3488
rect 201000 3476 201006 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 223868 3516 223896 3556
rect 235442 3544 235448 3556
rect 235500 3544 235506 3596
rect 241422 3544 241428 3596
rect 241480 3584 241486 3596
rect 244090 3584 244096 3596
rect 241480 3556 244096 3584
rect 241480 3544 241486 3556
rect 244090 3544 244096 3556
rect 244148 3544 244154 3596
rect 245470 3544 245476 3596
rect 245528 3584 245534 3596
rect 258046 3584 258074 3624
rect 262950 3612 262956 3624
rect 263008 3612 263014 3664
rect 264238 3612 264244 3664
rect 264296 3652 264302 3664
rect 264296 3624 266676 3652
rect 264296 3612 264302 3624
rect 245528 3556 258074 3584
rect 245528 3544 245534 3556
rect 261754 3544 261760 3596
rect 261812 3584 261818 3596
rect 262214 3584 262220 3596
rect 261812 3556 262220 3584
rect 261812 3544 261818 3556
rect 262214 3544 262220 3556
rect 262272 3544 262278 3596
rect 262858 3544 262864 3596
rect 262916 3584 262922 3596
rect 266538 3584 266544 3596
rect 262916 3556 266544 3584
rect 262916 3544 262922 3556
rect 266538 3544 266544 3556
rect 266596 3544 266602 3596
rect 266648 3584 266676 3624
rect 266722 3612 266728 3664
rect 266780 3652 266786 3664
rect 350442 3652 350448 3664
rect 266780 3624 350448 3652
rect 266780 3612 266786 3624
rect 350442 3612 350448 3624
rect 350500 3612 350506 3664
rect 356698 3612 356704 3664
rect 356756 3652 356762 3664
rect 369394 3652 369400 3664
rect 356756 3624 369400 3652
rect 356756 3612 356762 3624
rect 369394 3612 369400 3624
rect 369452 3612 369458 3664
rect 395338 3612 395344 3664
rect 395396 3652 395402 3664
rect 397730 3652 397736 3664
rect 395396 3624 397736 3652
rect 395396 3612 395402 3624
rect 397730 3612 397736 3624
rect 397788 3612 397794 3664
rect 399478 3612 399484 3664
rect 399536 3652 399542 3664
rect 450906 3652 450912 3664
rect 399536 3624 450912 3652
rect 399536 3612 399542 3624
rect 450906 3612 450912 3624
rect 450964 3612 450970 3664
rect 454678 3612 454684 3664
rect 454736 3652 454742 3664
rect 515950 3652 515956 3664
rect 454736 3624 515956 3652
rect 454736 3612 454742 3624
rect 515950 3612 515956 3624
rect 516008 3612 516014 3664
rect 527818 3652 527824 3664
rect 518866 3624 527824 3652
rect 273622 3584 273628 3596
rect 266648 3556 273628 3584
rect 273622 3544 273628 3556
rect 273680 3544 273686 3596
rect 293218 3544 293224 3596
rect 293276 3584 293282 3596
rect 294874 3584 294880 3596
rect 293276 3556 294880 3584
rect 293276 3544 293282 3556
rect 294874 3544 294880 3556
rect 294932 3544 294938 3596
rect 295978 3544 295984 3596
rect 296036 3584 296042 3596
rect 465166 3584 465172 3596
rect 296036 3556 465172 3584
rect 296036 3544 296042 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 469858 3584 469864 3596
rect 467156 3556 469864 3584
rect 467156 3544 467162 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 471238 3544 471244 3596
rect 471296 3584 471302 3596
rect 518866 3584 518894 3624
rect 527818 3612 527824 3624
rect 527876 3612 527882 3664
rect 471296 3556 518894 3584
rect 471296 3544 471302 3556
rect 520918 3544 520924 3596
rect 520976 3584 520982 3596
rect 523034 3584 523040 3596
rect 520976 3556 523040 3584
rect 520976 3544 520982 3556
rect 523034 3544 523040 3556
rect 523092 3544 523098 3596
rect 540238 3544 540244 3596
rect 540296 3584 540302 3596
rect 541986 3584 541992 3596
rect 540296 3556 541992 3584
rect 540296 3544 540302 3556
rect 541986 3544 541992 3556
rect 542044 3544 542050 3596
rect 547138 3544 547144 3596
rect 547196 3584 547202 3596
rect 552658 3584 552664 3596
rect 547196 3556 552664 3584
rect 547196 3544 547202 3556
rect 552658 3544 552664 3556
rect 552716 3544 552722 3596
rect 206244 3488 223896 3516
rect 206244 3476 206250 3488
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224862 3516 224868 3528
rect 224000 3488 224868 3516
rect 224000 3476 224006 3488
rect 224862 3476 224868 3488
rect 224920 3476 224926 3528
rect 230382 3476 230388 3528
rect 230440 3516 230446 3528
rect 231026 3516 231032 3528
rect 230440 3488 231032 3516
rect 230440 3476 230446 3488
rect 231026 3476 231032 3488
rect 231084 3476 231090 3528
rect 232222 3476 232228 3528
rect 232280 3516 232286 3528
rect 233142 3516 233148 3528
rect 232280 3488 233148 3516
rect 232280 3476 232286 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 245102 3476 245108 3528
rect 245160 3516 245166 3528
rect 270034 3516 270040 3528
rect 245160 3488 270040 3516
rect 245160 3476 245166 3488
rect 270034 3476 270040 3488
rect 270092 3476 270098 3528
rect 271138 3476 271144 3528
rect 271196 3516 271202 3528
rect 274818 3516 274824 3528
rect 271196 3488 274824 3516
rect 271196 3476 271202 3488
rect 274818 3476 274824 3488
rect 274876 3476 274882 3528
rect 276934 3476 276940 3528
rect 276992 3516 276998 3528
rect 449158 3516 449164 3528
rect 276992 3488 449164 3516
rect 276992 3476 276998 3488
rect 449158 3476 449164 3488
rect 449216 3476 449222 3528
rect 449268 3488 454034 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 200390 3448 200396 3460
rect 6512 3420 200396 3448
rect 6512 3408 6518 3420
rect 200390 3408 200396 3420
rect 200448 3408 200454 3460
rect 203886 3408 203892 3460
rect 203944 3448 203950 3460
rect 233602 3448 233608 3460
rect 203944 3420 233608 3448
rect 203944 3408 203950 3420
rect 233602 3408 233608 3420
rect 233660 3408 233666 3460
rect 234430 3408 234436 3460
rect 234488 3448 234494 3460
rect 237006 3448 237012 3460
rect 234488 3420 237012 3448
rect 234488 3408 234494 3420
rect 237006 3408 237012 3420
rect 237064 3408 237070 3460
rect 246574 3408 246580 3460
rect 246632 3448 246638 3460
rect 272426 3448 272432 3460
rect 246632 3420 272432 3448
rect 246632 3408 246638 3420
rect 272426 3408 272432 3420
rect 272484 3408 272490 3460
rect 282178 3408 282184 3460
rect 282236 3448 282242 3460
rect 283098 3448 283104 3460
rect 282236 3420 283104 3448
rect 282236 3408 282242 3420
rect 283098 3408 283104 3420
rect 283156 3408 283162 3460
rect 449268 3448 449296 3488
rect 287026 3420 449296 3448
rect 454006 3448 454034 3488
rect 457438 3476 457444 3528
rect 457496 3516 457502 3528
rect 534902 3516 534908 3528
rect 457496 3488 534908 3516
rect 457496 3476 457502 3488
rect 534902 3476 534908 3488
rect 534960 3476 534966 3528
rect 536098 3476 536104 3528
rect 536156 3516 536162 3528
rect 550266 3516 550272 3528
rect 536156 3488 550272 3516
rect 536156 3476 536162 3488
rect 550266 3476 550272 3488
rect 550324 3476 550330 3528
rect 479334 3448 479340 3460
rect 454006 3420 479340 3448
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 75178 3380 75184 3392
rect 66772 3352 75184 3380
rect 66772 3340 66778 3352
rect 75178 3340 75184 3352
rect 75236 3340 75242 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 86218 3380 86224 3392
rect 80940 3352 86224 3380
rect 80940 3340 80946 3352
rect 86218 3340 86224 3352
rect 86276 3340 86282 3392
rect 110506 3340 110512 3392
rect 110564 3380 110570 3392
rect 111702 3380 111708 3392
rect 110564 3352 111708 3380
rect 110564 3340 110570 3352
rect 111702 3340 111708 3352
rect 111760 3340 111766 3392
rect 141234 3340 141240 3392
rect 141292 3380 141298 3392
rect 142062 3380 142068 3392
rect 141292 3352 142068 3380
rect 141292 3340 141298 3352
rect 142062 3340 142068 3352
rect 142120 3340 142126 3392
rect 150618 3340 150624 3392
rect 150676 3380 150682 3392
rect 225230 3380 225236 3392
rect 150676 3352 225236 3380
rect 150676 3340 150682 3352
rect 225230 3340 225236 3352
rect 225288 3340 225294 3392
rect 242710 3340 242716 3392
rect 242768 3380 242774 3392
rect 242768 3352 248414 3380
rect 242768 3340 242774 3352
rect 59630 3272 59636 3324
rect 59688 3312 59694 3324
rect 68278 3312 68284 3324
rect 59688 3284 68284 3312
rect 59688 3272 59694 3284
rect 68278 3272 68284 3284
rect 68336 3272 68342 3324
rect 169570 3272 169576 3324
rect 169628 3312 169634 3324
rect 170398 3312 170404 3324
rect 169628 3284 170404 3312
rect 169628 3272 169634 3284
rect 170398 3272 170404 3284
rect 170456 3272 170462 3324
rect 205082 3272 205088 3324
rect 205140 3312 205146 3324
rect 217318 3312 217324 3324
rect 205140 3284 217324 3312
rect 205140 3272 205146 3284
rect 217318 3272 217324 3284
rect 217376 3272 217382 3324
rect 242434 3272 242440 3324
rect 242492 3312 242498 3324
rect 246390 3312 246396 3324
rect 242492 3284 246396 3312
rect 242492 3272 242498 3284
rect 246390 3272 246396 3284
rect 246448 3272 246454 3324
rect 248386 3312 248414 3352
rect 280982 3340 280988 3392
rect 281040 3380 281046 3392
rect 287026 3380 287054 3420
rect 479334 3408 479340 3420
rect 479392 3408 479398 3460
rect 486418 3408 486424 3460
rect 486476 3448 486482 3460
rect 488810 3448 488816 3460
rect 486476 3420 488816 3448
rect 486476 3408 486482 3420
rect 488810 3408 488816 3420
rect 488868 3408 488874 3460
rect 547874 3448 547880 3460
rect 489886 3420 547880 3448
rect 281040 3352 287054 3380
rect 281040 3340 281046 3352
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 311250 3340 311256 3392
rect 311308 3380 311314 3392
rect 312630 3380 312636 3392
rect 311308 3352 312636 3380
rect 311308 3340 311314 3352
rect 312630 3340 312636 3352
rect 312688 3340 312694 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 318150 3340 318156 3392
rect 318208 3380 318214 3392
rect 319714 3380 319720 3392
rect 318208 3352 319720 3380
rect 318208 3340 318214 3352
rect 319714 3340 319720 3352
rect 319772 3340 319778 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 331858 3340 331864 3392
rect 331916 3380 331922 3392
rect 332686 3380 332692 3392
rect 331916 3352 332692 3380
rect 331916 3340 331922 3352
rect 332686 3340 332692 3352
rect 332744 3340 332750 3392
rect 335998 3340 336004 3392
rect 336056 3380 336062 3392
rect 337470 3380 337476 3392
rect 336056 3352 337476 3380
rect 336056 3340 336062 3352
rect 337470 3340 337476 3352
rect 337528 3340 337534 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 342990 3340 342996 3392
rect 343048 3380 343054 3392
rect 344554 3380 344560 3392
rect 343048 3352 344560 3380
rect 343048 3340 343054 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 345658 3340 345664 3392
rect 345716 3380 345722 3392
rect 348050 3380 348056 3392
rect 345716 3352 348056 3380
rect 345716 3340 345722 3352
rect 348050 3340 348056 3352
rect 348108 3340 348114 3392
rect 360838 3340 360844 3392
rect 360896 3380 360902 3392
rect 363506 3380 363512 3392
rect 360896 3352 363512 3380
rect 360896 3340 360902 3352
rect 363506 3340 363512 3352
rect 363564 3340 363570 3392
rect 367830 3340 367836 3392
rect 367888 3380 367894 3392
rect 370590 3380 370596 3392
rect 367888 3352 370596 3380
rect 367888 3340 367894 3352
rect 370590 3340 370596 3352
rect 370648 3340 370654 3392
rect 374638 3340 374644 3392
rect 374696 3380 374702 3392
rect 377674 3380 377680 3392
rect 374696 3352 377680 3380
rect 374696 3340 374702 3352
rect 377674 3340 377680 3352
rect 377732 3340 377738 3392
rect 378778 3340 378784 3392
rect 378836 3380 378842 3392
rect 381170 3380 381176 3392
rect 378836 3352 381176 3380
rect 378836 3340 378842 3352
rect 381170 3340 381176 3352
rect 381228 3340 381234 3392
rect 382918 3340 382924 3392
rect 382976 3380 382982 3392
rect 384758 3380 384764 3392
rect 382976 3352 384764 3380
rect 382976 3340 382982 3352
rect 384758 3340 384764 3352
rect 384816 3340 384822 3392
rect 389818 3340 389824 3392
rect 389876 3380 389882 3392
rect 391842 3380 391848 3392
rect 389876 3352 391848 3380
rect 389876 3340 389882 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 403618 3340 403624 3392
rect 403676 3380 403682 3392
rect 408402 3380 408408 3392
rect 403676 3352 408408 3380
rect 403676 3340 403682 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 421374 3380 421380 3392
rect 414716 3352 421380 3380
rect 414716 3340 414722 3352
rect 421374 3340 421380 3352
rect 421432 3340 421438 3392
rect 421558 3340 421564 3392
rect 421616 3380 421622 3392
rect 427262 3380 427268 3392
rect 421616 3352 427268 3380
rect 421616 3340 421622 3352
rect 427262 3340 427268 3352
rect 427320 3340 427326 3392
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 442258 3340 442264 3392
rect 442316 3380 442322 3392
rect 446214 3380 446220 3392
rect 442316 3352 446220 3380
rect 442316 3340 442322 3352
rect 446214 3340 446220 3352
rect 446272 3340 446278 3392
rect 449158 3340 449164 3392
rect 449216 3380 449222 3392
rect 449216 3352 456794 3380
rect 449216 3340 449222 3352
rect 248782 3312 248788 3324
rect 248386 3284 248788 3312
rect 248782 3272 248788 3284
rect 248840 3272 248846 3324
rect 324958 3272 324964 3324
rect 325016 3312 325022 3324
rect 326798 3312 326804 3324
rect 325016 3284 326804 3312
rect 325016 3272 325022 3284
rect 326798 3272 326804 3284
rect 326856 3272 326862 3324
rect 31294 3204 31300 3256
rect 31352 3244 31358 3256
rect 33778 3244 33784 3256
rect 31352 3216 33784 3244
rect 31352 3204 31358 3216
rect 33778 3204 33784 3216
rect 33836 3204 33842 3256
rect 143534 3204 143540 3256
rect 143592 3244 143598 3256
rect 144822 3244 144828 3256
rect 143592 3216 144828 3244
rect 143592 3204 143598 3216
rect 144822 3204 144828 3216
rect 144880 3204 144886 3256
rect 168374 3204 168380 3256
rect 168432 3244 168438 3256
rect 169662 3244 169668 3256
rect 168432 3216 169668 3244
rect 168432 3204 168438 3216
rect 169662 3204 169668 3216
rect 169720 3204 169726 3256
rect 173158 3204 173164 3256
rect 173216 3244 173222 3256
rect 174538 3244 174544 3256
rect 173216 3216 174544 3244
rect 173216 3204 173222 3216
rect 174538 3204 174544 3216
rect 174596 3204 174602 3256
rect 222746 3204 222752 3256
rect 222804 3244 222810 3256
rect 229738 3244 229744 3256
rect 222804 3216 229744 3244
rect 222804 3204 222810 3216
rect 229738 3204 229744 3216
rect 229796 3204 229802 3256
rect 242158 3204 242164 3256
rect 242216 3244 242222 3256
rect 245194 3244 245200 3256
rect 242216 3216 245200 3244
rect 242216 3204 242222 3216
rect 245194 3204 245200 3216
rect 245252 3204 245258 3256
rect 250438 3204 250444 3256
rect 250496 3244 250502 3256
rect 254670 3244 254676 3256
rect 250496 3216 254676 3244
rect 250496 3204 250502 3216
rect 254670 3204 254676 3216
rect 254728 3204 254734 3256
rect 385678 3204 385684 3256
rect 385736 3244 385742 3256
rect 387150 3244 387156 3256
rect 385736 3216 387156 3244
rect 385736 3204 385742 3216
rect 387150 3204 387156 3216
rect 387208 3204 387214 3256
rect 456766 3244 456794 3352
rect 485038 3340 485044 3392
rect 485096 3380 485102 3392
rect 489886 3380 489914 3420
rect 547874 3408 547880 3420
rect 547932 3408 547938 3460
rect 558178 3408 558184 3460
rect 558236 3448 558242 3460
rect 565630 3448 565636 3460
rect 558236 3420 565636 3448
rect 558236 3408 558242 3420
rect 565630 3408 565636 3420
rect 565688 3408 565694 3460
rect 485096 3352 489914 3380
rect 485096 3340 485102 3352
rect 490558 3340 490564 3392
rect 490616 3380 490622 3392
rect 492306 3380 492312 3392
rect 490616 3352 492312 3380
rect 490616 3340 490622 3352
rect 492306 3340 492312 3352
rect 492364 3340 492370 3392
rect 497458 3340 497464 3392
rect 497516 3380 497522 3392
rect 499390 3380 499396 3392
rect 497516 3352 499396 3380
rect 497516 3340 497522 3352
rect 499390 3340 499396 3352
rect 499448 3340 499454 3392
rect 515398 3340 515404 3392
rect 515456 3380 515462 3392
rect 517146 3380 517152 3392
rect 515456 3352 517152 3380
rect 515456 3340 515462 3352
rect 517146 3340 517152 3352
rect 517204 3340 517210 3392
rect 465718 3272 465724 3324
rect 465776 3312 465782 3324
rect 467466 3312 467472 3324
rect 465776 3284 467472 3312
rect 465776 3272 465782 3284
rect 467466 3272 467472 3284
rect 467524 3272 467530 3324
rect 482278 3272 482284 3324
rect 482336 3312 482342 3324
rect 486418 3312 486424 3324
rect 482336 3284 486424 3312
rect 482336 3272 482342 3284
rect 486418 3272 486424 3284
rect 486476 3272 486482 3324
rect 500310 3272 500316 3324
rect 500368 3312 500374 3324
rect 502978 3312 502984 3324
rect 500368 3284 502984 3312
rect 500368 3272 500374 3284
rect 502978 3272 502984 3284
rect 503036 3272 503042 3324
rect 580258 3272 580264 3324
rect 580316 3312 580322 3324
rect 580994 3312 581000 3324
rect 580316 3284 581000 3312
rect 580316 3272 580322 3284
rect 580994 3272 581000 3284
rect 581052 3272 581058 3324
rect 458082 3244 458088 3256
rect 456766 3216 458088 3244
rect 458082 3204 458088 3216
rect 458140 3204 458146 3256
rect 48958 3136 48964 3188
rect 49016 3176 49022 3188
rect 53098 3176 53104 3188
rect 49016 3148 53104 3176
rect 49016 3136 49022 3148
rect 53098 3136 53104 3148
rect 53156 3136 53162 3188
rect 235810 3136 235816 3188
rect 235868 3176 235874 3188
rect 238018 3176 238024 3188
rect 235868 3148 238024 3176
rect 235868 3136 235874 3148
rect 238018 3136 238024 3148
rect 238076 3136 238082 3188
rect 239306 3136 239312 3188
rect 239364 3176 239370 3188
rect 240778 3176 240784 3188
rect 239364 3148 240784 3176
rect 239364 3136 239370 3148
rect 240778 3136 240784 3148
rect 240836 3136 240842 3188
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 201954 3108 201960 3120
rect 15988 3080 201960 3108
rect 15988 3068 15994 3080
rect 201954 3068 201960 3080
rect 202012 3068 202018 3120
rect 242526 3068 242532 3120
rect 242584 3108 242590 3120
rect 247586 3108 247592 3120
rect 242584 3080 247592 3108
rect 242584 3068 242590 3080
rect 247586 3068 247592 3080
rect 247644 3068 247650 3120
rect 413278 3068 413284 3120
rect 413336 3108 413342 3120
rect 420178 3108 420184 3120
rect 413336 3080 420184 3108
rect 413336 3068 413342 3080
rect 420178 3068 420184 3080
rect 420236 3068 420242 3120
rect 542998 3068 543004 3120
rect 543056 3108 543062 3120
rect 545482 3108 545488 3120
rect 543056 3080 545488 3108
rect 543056 3068 543062 3080
rect 545482 3068 545488 3080
rect 545540 3068 545546 3120
rect 554038 3068 554044 3120
rect 554096 3108 554102 3120
rect 556154 3108 556160 3120
rect 554096 3080 556160 3108
rect 554096 3068 554102 3080
rect 556154 3068 556160 3080
rect 556212 3068 556218 3120
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 14458 3040 14464 3052
rect 8812 3012 14464 3040
rect 8812 3000 8818 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 104526 3000 104532 3052
rect 104584 3040 104590 3052
rect 105538 3040 105544 3052
rect 104584 3012 105544 3040
rect 104584 3000 104590 3012
rect 105538 3000 105544 3012
rect 105596 3000 105602 3052
rect 184934 3000 184940 3052
rect 184992 3040 184998 3052
rect 187050 3040 187056 3052
rect 184992 3012 187056 3040
rect 184992 3000 184998 3012
rect 187050 3000 187056 3012
rect 187108 3000 187114 3052
rect 233418 3000 233424 3052
rect 233476 3040 233482 3052
rect 234522 3040 234528 3052
rect 233476 3012 234528 3040
rect 233476 3000 233482 3012
rect 234522 3000 234528 3012
rect 234580 3000 234586 3052
rect 364978 3000 364984 3052
rect 365036 3040 365042 3052
rect 367002 3040 367008 3052
rect 365036 3012 367008 3040
rect 365036 3000 365042 3012
rect 367002 3000 367008 3012
rect 367060 3000 367066 3052
rect 369118 3000 369124 3052
rect 369176 3040 369182 3052
rect 371694 3040 371700 3052
rect 369176 3012 371700 3040
rect 369176 3000 369182 3012
rect 371694 3000 371700 3012
rect 371752 3000 371758 3052
rect 377398 3000 377404 3052
rect 377456 3040 377462 3052
rect 379974 3040 379980 3052
rect 377456 3012 379980 3040
rect 377456 3000 377462 3012
rect 379974 3000 379980 3012
rect 380032 3000 380038 3052
rect 435358 3000 435364 3052
rect 435416 3040 435422 3052
rect 437934 3040 437940 3052
rect 435416 3012 437940 3040
rect 435416 3000 435422 3012
rect 437934 3000 437940 3012
rect 437992 3000 437998 3052
rect 504358 3000 504364 3052
rect 504416 3040 504422 3052
rect 510062 3040 510068 3052
rect 504416 3012 510068 3040
rect 504416 3000 504422 3012
rect 510062 3000 510068 3012
rect 510120 3000 510126 3052
rect 511258 3000 511264 3052
rect 511316 3040 511322 3052
rect 513558 3040 513564 3052
rect 511316 3012 513564 3040
rect 511316 3000 511322 3012
rect 513558 3000 513564 3012
rect 513616 3000 513622 3052
rect 529198 3000 529204 3052
rect 529256 3040 529262 3052
rect 531314 3040 531320 3052
rect 529256 3012 531320 3040
rect 529256 3000 529262 3012
rect 531314 3000 531320 3012
rect 531372 3000 531378 3052
rect 312538 2932 312544 2984
rect 312596 2972 312602 2984
rect 315022 2972 315028 2984
rect 312596 2944 315028 2972
rect 312596 2932 312602 2944
rect 315022 2932 315028 2944
rect 315080 2932 315086 2984
rect 446398 2932 446404 2984
rect 446456 2972 446462 2984
rect 452102 2972 452108 2984
rect 446456 2944 452108 2972
rect 446456 2932 446462 2944
rect 452102 2932 452108 2944
rect 452160 2932 452166 2984
rect 493318 2932 493324 2984
rect 493376 2972 493382 2984
rect 495894 2972 495900 2984
rect 493376 2944 495900 2972
rect 493376 2932 493382 2944
rect 495894 2932 495900 2944
rect 495952 2932 495958 2984
rect 522298 2932 522304 2984
rect 522356 2972 522362 2984
rect 524230 2972 524236 2984
rect 522356 2944 524236 2972
rect 522356 2932 522362 2944
rect 524230 2932 524236 2944
rect 524288 2932 524294 2984
rect 530670 2932 530676 2984
rect 530728 2972 530734 2984
rect 532510 2972 532516 2984
rect 530728 2944 532516 2972
rect 530728 2932 530734 2944
rect 532510 2932 532516 2944
rect 532568 2932 532574 2984
rect 275278 2864 275284 2916
rect 275336 2904 275342 2916
rect 279510 2904 279516 2916
rect 275336 2876 279516 2904
rect 275336 2864 275342 2876
rect 279510 2864 279516 2876
rect 279568 2864 279574 2916
rect 472710 2864 472716 2916
rect 472768 2904 472774 2916
rect 474550 2904 474556 2916
rect 472768 2876 474556 2904
rect 472768 2864 472774 2876
rect 474550 2864 474556 2876
rect 474608 2864 474614 2916
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 202788 700952 202840 701004
rect 251180 700952 251232 701004
rect 248328 700884 248380 700936
rect 348792 700884 348844 700936
rect 154120 700816 154172 700868
rect 255320 700816 255372 700868
rect 137836 700748 137888 700800
rect 253940 700748 253992 700800
rect 245568 700680 245620 700732
rect 413652 700680 413704 700732
rect 89168 700612 89220 700664
rect 256792 700612 256844 700664
rect 72976 700544 73028 700596
rect 256700 700544 256752 700596
rect 40500 700476 40552 700528
rect 41328 700476 41380 700528
rect 242808 700476 242860 700528
rect 478512 700476 478564 700528
rect 24308 700408 24360 700460
rect 259552 700408 259604 700460
rect 8116 700340 8168 700392
rect 259460 700340 259512 700392
rect 295984 700340 296036 700392
rect 300124 700340 300176 700392
rect 241336 700272 241388 700324
rect 543464 700272 543516 700324
rect 218980 700204 219032 700256
rect 252560 700204 252612 700256
rect 251088 700136 251140 700188
rect 283840 700136 283892 700188
rect 249708 700068 249760 700120
rect 267648 700068 267700 700120
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 233148 699660 233200 699712
rect 235172 699660 235224 699712
rect 359464 699660 359516 699712
rect 364984 699660 365036 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 461584 699660 461636 699712
rect 462320 699660 462372 699712
rect 526444 699660 526496 699712
rect 527180 699660 527232 699712
rect 237288 696940 237340 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 260840 683204 260892 683256
rect 238576 683136 238628 683188
rect 580172 683136 580224 683188
rect 3424 670760 3476 670812
rect 262220 670760 262272 670812
rect 235908 670692 235960 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 262312 656888 262364 656940
rect 234528 643084 234580 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 263600 632068 263652 632120
rect 235816 630640 235868 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 264980 618264 265032 618316
rect 234436 616836 234488 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 263692 605820 263744 605872
rect 231676 590656 231728 590708
rect 579804 590656 579856 590708
rect 371700 585352 371752 585404
rect 513564 585352 513616 585404
rect 446404 585284 446456 585336
rect 513380 585284 513432 585336
rect 425704 585216 425756 585268
rect 516416 585216 516468 585268
rect 489184 584468 489236 584520
rect 513932 584468 513984 584520
rect 485044 584400 485096 584452
rect 513564 584400 513616 584452
rect 371792 584332 371844 584384
rect 513748 584332 513800 584384
rect 500224 584264 500276 584316
rect 516324 584264 516376 584316
rect 493324 584196 493376 584248
rect 513840 584196 513892 584248
rect 490564 584128 490616 584180
rect 513656 584128 513708 584180
rect 483664 584060 483716 584112
rect 513380 584060 513432 584112
rect 430580 583992 430632 584044
rect 516232 583992 516284 584044
rect 427820 583924 427872 583976
rect 513288 583924 513340 583976
rect 444748 583856 444800 583908
rect 447784 583856 447836 583908
rect 497464 583856 497516 583908
rect 513472 583856 513524 583908
rect 516140 583720 516192 583772
rect 524420 583720 524472 583772
rect 371608 581068 371660 581120
rect 374000 581068 374052 581120
rect 371332 581000 371384 581052
rect 378232 581000 378284 581052
rect 378784 580252 378836 580304
rect 427820 580252 427872 580304
rect 371516 579776 371568 579828
rect 377036 579776 377088 579828
rect 371608 579708 371660 579760
rect 378784 579708 378836 579760
rect 3332 579640 3384 579692
rect 266360 579640 266412 579692
rect 371700 579640 371752 579692
rect 380164 579640 380216 579692
rect 444748 579640 444800 579692
rect 447876 579640 447928 579692
rect 444932 578416 444984 578468
rect 448152 578416 448204 578468
rect 371332 578280 371384 578332
rect 375472 578280 375524 578332
rect 371700 578212 371752 578264
rect 379152 578212 379204 578264
rect 371240 578076 371292 578128
rect 371792 578076 371844 578128
rect 378140 577464 378192 577516
rect 430580 577464 430632 577516
rect 371424 576988 371476 577040
rect 376760 576988 376812 577040
rect 371608 576920 371660 576972
rect 378140 576920 378192 576972
rect 371700 576852 371752 576904
rect 379060 576852 379112 576904
rect 371608 576104 371660 576156
rect 425704 576104 425756 576156
rect 371700 575492 371752 575544
rect 376944 575492 376996 575544
rect 444748 575492 444800 575544
rect 448244 575492 448296 575544
rect 444564 574064 444616 574116
rect 447968 574064 448020 574116
rect 371608 571480 371660 571532
rect 375380 571480 375432 571532
rect 444840 571480 444892 571532
rect 448060 571480 448112 571532
rect 371516 570256 371568 570308
rect 376208 570256 376260 570308
rect 371608 569984 371660 570036
rect 376024 569984 376076 570036
rect 371700 569916 371752 569968
rect 376852 569916 376904 569968
rect 516140 568896 516192 568948
rect 520372 568896 520424 568948
rect 444932 568556 444984 568608
rect 449164 568556 449216 568608
rect 516232 568556 516284 568608
rect 524604 568556 524656 568608
rect 516508 568012 516560 568064
rect 516784 568012 516836 568064
rect 371516 567876 371568 567928
rect 372988 567876 373040 567928
rect 371516 567740 371568 567792
rect 371700 567740 371752 567792
rect 371608 567672 371660 567724
rect 374644 567672 374696 567724
rect 516232 567332 516284 567384
rect 521752 567332 521804 567384
rect 516140 567264 516192 567316
rect 519360 567264 519412 567316
rect 516232 567196 516284 567248
rect 516876 567196 516928 567248
rect 516600 567128 516652 567180
rect 516876 567060 516928 567112
rect 516508 566992 516560 567044
rect 516784 566992 516836 567044
rect 371792 566176 371844 566228
rect 374184 566176 374236 566228
rect 516508 566040 516560 566092
rect 520464 566040 520516 566092
rect 3424 565836 3476 565888
rect 267740 565836 267792 565888
rect 371792 565836 371844 565888
rect 373264 565836 373316 565888
rect 516416 565836 516468 565888
rect 521936 565836 521988 565888
rect 371792 564680 371844 564732
rect 374276 564680 374328 564732
rect 516508 564680 516560 564732
rect 520556 564680 520608 564732
rect 444380 564544 444432 564596
rect 446496 564544 446548 564596
rect 516416 564476 516468 564528
rect 519268 564476 519320 564528
rect 516324 563728 516376 563780
rect 520280 563728 520332 563780
rect 516324 563252 516376 563304
rect 518992 563252 519044 563304
rect 371792 563048 371844 563100
rect 374368 563048 374420 563100
rect 445668 563048 445720 563100
rect 450544 563048 450596 563100
rect 516324 563048 516376 563100
rect 517796 563048 517848 563100
rect 371792 562504 371844 562556
rect 374460 562504 374512 562556
rect 516324 562504 516376 562556
rect 519084 562504 519136 562556
rect 516324 561960 516376 562012
rect 517888 561960 517940 562012
rect 516324 561416 516376 561468
rect 517980 561416 518032 561468
rect 444380 561144 444432 561196
rect 446588 561144 446640 561196
rect 371792 560872 371844 560924
rect 375564 560872 375616 560924
rect 371792 560328 371844 560380
rect 376116 560328 376168 560380
rect 371792 559104 371844 559156
rect 374552 559104 374604 559156
rect 516324 558968 516376 559020
rect 524696 558968 524748 559020
rect 371884 558900 371936 558952
rect 377128 558900 377180 558952
rect 516508 558900 516560 558952
rect 525800 558900 525852 558952
rect 371792 558152 371844 558204
rect 374092 558152 374144 558204
rect 371792 558016 371844 558068
rect 375656 558016 375708 558068
rect 441620 558016 441672 558068
rect 516508 557744 516560 557796
rect 519176 557744 519228 557796
rect 516324 557676 516376 557728
rect 523040 557676 523092 557728
rect 444380 557608 444432 557660
rect 447140 557608 447192 557660
rect 516784 557608 516836 557660
rect 517060 557608 517112 557660
rect 521844 557608 521896 557660
rect 516600 557540 516652 557592
rect 502984 557064 503036 557116
rect 516140 557064 516192 557116
rect 501604 556996 501656 557048
rect 516324 556996 516376 557048
rect 486424 556928 486476 556980
rect 516600 556928 516652 556980
rect 454684 556860 454736 556912
rect 516416 556860 516468 556912
rect 370504 556792 370556 556844
rect 441712 556792 441764 556844
rect 513380 556792 513432 556844
rect 371792 556248 371844 556300
rect 372896 556248 372948 556300
rect 516140 556248 516192 556300
rect 521660 556248 521712 556300
rect 516232 556180 516284 556232
rect 524512 556180 524564 556232
rect 376024 556112 376076 556164
rect 516876 556112 516928 556164
rect 373264 556044 373316 556096
rect 441620 556044 441672 556096
rect 376116 555976 376168 556028
rect 444472 555976 444524 556028
rect 503352 555908 503404 555960
rect 513472 555908 513524 555960
rect 503260 555840 503312 555892
rect 513564 555840 513616 555892
rect 503168 555772 503220 555824
rect 513656 555772 513708 555824
rect 503076 555704 503128 555756
rect 513748 555704 513800 555756
rect 482284 555636 482336 555688
rect 516508 555636 516560 555688
rect 464344 555568 464396 555620
rect 516968 555568 517020 555620
rect 456708 555500 456760 555552
rect 513840 555500 513892 555552
rect 449256 555432 449308 555484
rect 516692 555432 516744 555484
rect 516784 554752 516836 554804
rect 517520 554752 517572 554804
rect 435180 554684 435232 554736
rect 506848 554684 506900 554736
rect 198648 554140 198700 554192
rect 366916 554140 366968 554192
rect 302884 554072 302936 554124
rect 510896 554072 510948 554124
rect 198556 554004 198608 554056
rect 438952 554004 439004 554056
rect 3424 553392 3476 553444
rect 266452 553392 266504 553444
rect 512920 553392 512972 553444
rect 514760 553392 514812 553444
rect 368940 551896 368992 551948
rect 369308 551896 369360 551948
rect 448152 541628 448204 541680
rect 521936 541628 521988 541680
rect 230388 536800 230440 536852
rect 580172 536800 580224 536852
rect 448244 536052 448296 536104
rect 520556 536052 520608 536104
rect 3424 527144 3476 527196
rect 267832 527144 267884 527196
rect 449164 526396 449216 526448
rect 449348 526396 449400 526448
rect 517888 526396 517940 526448
rect 230296 524424 230348 524476
rect 580172 524424 580224 524476
rect 446496 523676 446548 523728
rect 525800 523676 525852 523728
rect 376208 522928 376260 522980
rect 376668 522928 376720 522980
rect 450544 522316 450596 522368
rect 524696 522316 524748 522368
rect 376668 522248 376720 522300
rect 454040 522248 454092 522300
rect 454684 522248 454736 522300
rect 448060 520888 448112 520940
rect 517796 520888 517848 520940
rect 447876 517828 447928 517880
rect 448428 517828 448480 517880
rect 448428 517488 448480 517540
rect 516416 517488 516468 517540
rect 520464 517488 520516 517540
rect 369124 516944 369176 516996
rect 369492 516944 369544 516996
rect 516140 516060 516192 516112
rect 519268 516060 519320 516112
rect 3424 514768 3476 514820
rect 270500 514768 270552 514820
rect 447876 514768 447928 514820
rect 516140 514768 516192 514820
rect 507860 514020 507912 514072
rect 513380 514020 513432 514072
rect 517152 514020 517204 514072
rect 518164 514020 518216 514072
rect 524604 514020 524656 514072
rect 444380 513748 444432 513800
rect 444932 513748 444984 513800
rect 446404 513748 446456 513800
rect 444564 512728 444616 512780
rect 483664 512728 483716 512780
rect 516140 512728 516192 512780
rect 520372 512728 520424 512780
rect 447784 512660 447836 512712
rect 513748 512660 513800 512712
rect 445392 512592 445444 512644
rect 514852 512592 514904 512644
rect 445668 511912 445720 511964
rect 485044 511912 485096 511964
rect 369124 511776 369176 511828
rect 369400 511776 369452 511828
rect 370964 511164 371016 511216
rect 372988 511164 373040 511216
rect 517704 510620 517756 510672
rect 518900 510620 518952 510672
rect 370964 510008 371016 510060
rect 374644 510008 374696 510060
rect 374920 510008 374972 510060
rect 445668 509940 445720 509992
rect 452660 509940 452712 509992
rect 489184 509940 489236 509992
rect 445576 509872 445628 509924
rect 451280 509872 451332 509924
rect 490564 509872 490616 509924
rect 516140 509872 516192 509924
rect 521752 509872 521804 509924
rect 516140 508784 516192 508836
rect 519360 508784 519412 508836
rect 445668 508512 445720 508564
rect 450176 508512 450228 508564
rect 493324 508512 493376 508564
rect 445576 507832 445628 507884
rect 519360 507832 519412 507884
rect 520648 507832 520700 507884
rect 449164 507764 449216 507816
rect 503352 507764 503404 507816
rect 516140 507764 516192 507816
rect 521936 507764 521988 507816
rect 445576 507152 445628 507204
rect 450084 507152 450136 507204
rect 497464 507152 497516 507204
rect 445668 507084 445720 507136
rect 449992 507084 450044 507136
rect 500224 507084 500276 507136
rect 370964 506472 371016 506524
rect 374184 506472 374236 506524
rect 374828 506472 374880 506524
rect 445576 505860 445628 505912
rect 448520 505860 448572 505912
rect 449256 505860 449308 505912
rect 369124 505520 369176 505572
rect 369492 505520 369544 505572
rect 370044 505452 370096 505504
rect 373264 505452 373316 505504
rect 516968 505384 517020 505436
rect 517612 505384 517664 505436
rect 520372 505384 520424 505436
rect 445668 505112 445720 505164
rect 449900 505112 449952 505164
rect 448428 505044 448480 505096
rect 452752 505044 452804 505096
rect 449900 504976 449952 505028
rect 450544 504976 450596 505028
rect 503260 505044 503312 505096
rect 516140 505044 516192 505096
rect 520556 505044 520608 505096
rect 458180 504432 458232 504484
rect 464344 504432 464396 504484
rect 445668 504364 445720 504416
rect 448612 504364 448664 504416
rect 501604 504364 501656 504416
rect 370964 504160 371016 504212
rect 372620 504160 372672 504212
rect 373080 504160 373132 504212
rect 445300 503684 445352 503736
rect 458180 503684 458232 503736
rect 458824 503684 458876 503736
rect 446404 503616 446456 503668
rect 447876 503616 447928 503668
rect 370964 503140 371016 503192
rect 374276 503140 374328 503192
rect 445208 502256 445260 502308
rect 503168 502256 503220 502308
rect 459560 501576 459612 501628
rect 460204 501576 460256 501628
rect 486424 501576 486476 501628
rect 516876 501372 516928 501424
rect 518256 501372 518308 501424
rect 520280 501372 520332 501424
rect 3056 500964 3108 501016
rect 269120 500964 269172 501016
rect 445300 500964 445352 501016
rect 459560 500964 459612 501016
rect 445484 500896 445536 500948
rect 503076 500896 503128 500948
rect 445576 500828 445628 500880
rect 482284 500828 482336 500880
rect 445668 500760 445720 500812
rect 456708 500760 456760 500812
rect 516140 500760 516192 500812
rect 518992 500760 519044 500812
rect 516140 500488 516192 500540
rect 517796 500488 517848 500540
rect 456708 500352 456760 500404
rect 457444 500352 457496 500404
rect 372712 500284 372764 500336
rect 373264 500284 373316 500336
rect 370964 499604 371016 499656
rect 374368 499604 374420 499656
rect 444656 499468 444708 499520
rect 454040 499468 454092 499520
rect 466828 498788 466880 498840
rect 467748 498788 467800 498840
rect 502984 498788 503036 498840
rect 370964 498448 371016 498500
rect 374460 498448 374512 498500
rect 516140 498448 516192 498500
rect 519084 498448 519136 498500
rect 445576 498176 445628 498228
rect 466828 498176 466880 498228
rect 516140 498108 516192 498160
rect 517888 498108 517940 498160
rect 445484 497768 445536 497820
rect 449256 497768 449308 497820
rect 445576 496952 445628 497004
rect 447508 496952 447560 497004
rect 445760 496816 445812 496868
rect 446312 496816 446364 496868
rect 447140 496816 447192 496868
rect 449348 496816 449400 496868
rect 516232 495456 516284 495508
rect 517520 495456 517572 495508
rect 517980 495456 518032 495508
rect 370964 494776 371016 494828
rect 375564 494776 375616 494828
rect 376208 494776 376260 494828
rect 445300 494708 445352 494760
rect 445576 494708 445628 494760
rect 445300 494572 445352 494624
rect 446128 494572 446180 494624
rect 448152 494572 448204 494624
rect 442448 494028 442500 494080
rect 442908 494028 442960 494080
rect 452752 494028 452804 494080
rect 370964 493960 371016 494012
rect 375564 493960 375616 494012
rect 376116 493960 376168 494012
rect 446220 493960 446272 494012
rect 448244 493960 448296 494012
rect 516232 493960 516284 494012
rect 525800 493960 525852 494012
rect 445300 493348 445352 493400
rect 446220 493348 446272 493400
rect 370780 493280 370832 493332
rect 377128 493280 377180 493332
rect 444656 493280 444708 493332
rect 446404 493280 446456 493332
rect 446956 493280 447008 493332
rect 516140 492600 516192 492652
rect 524696 492600 524748 492652
rect 370872 492328 370924 492380
rect 374552 492328 374604 492380
rect 377220 492328 377272 492380
rect 448796 491648 448848 491700
rect 450636 491648 450688 491700
rect 369124 491308 369176 491360
rect 369308 491308 369360 491360
rect 443552 491308 443604 491360
rect 445944 491240 445996 491292
rect 443920 491172 443972 491224
rect 447140 491172 447192 491224
rect 516140 491172 516192 491224
rect 519176 491172 519228 491224
rect 522120 491172 522172 491224
rect 445300 491036 445352 491088
rect 445944 491036 445996 491088
rect 448060 491036 448112 491088
rect 370964 490288 371016 490340
rect 374092 490288 374144 490340
rect 374552 490288 374604 490340
rect 516692 489812 516744 489864
rect 521844 489812 521896 489864
rect 370412 489336 370464 489388
rect 370688 489336 370740 489388
rect 443092 488724 443144 488776
rect 447416 488724 447468 488776
rect 441896 488520 441948 488572
rect 442356 488520 442408 488572
rect 517244 488452 517296 488504
rect 523040 488452 523092 488504
rect 369400 488044 369452 488096
rect 369768 488044 369820 488096
rect 375656 488044 375708 488096
rect 444656 487840 444708 487892
rect 446496 487840 446548 487892
rect 445300 487296 445352 487348
rect 448796 487296 448848 487348
rect 445484 487160 445536 487212
rect 448704 487160 448756 487212
rect 516140 486412 516192 486464
rect 520924 486412 520976 486464
rect 524512 486412 524564 486464
rect 446588 486004 446640 486056
rect 513472 486004 513524 486056
rect 445484 485800 445536 485852
rect 445852 485800 445904 485852
rect 446588 485800 446640 485852
rect 445116 485732 445168 485784
rect 513380 485732 513432 485784
rect 516140 485732 516192 485784
rect 521660 485732 521712 485784
rect 370964 485256 371016 485308
rect 372896 485256 372948 485308
rect 447324 485052 447376 485104
rect 513748 485052 513800 485104
rect 369124 484848 369176 484900
rect 369124 484644 369176 484696
rect 445484 484576 445536 484628
rect 447324 484576 447376 484628
rect 448704 484304 448756 484356
rect 449348 484304 449400 484356
rect 516232 484304 516284 484356
rect 513104 484236 513156 484288
rect 514760 484236 514812 484288
rect 444656 484168 444708 484220
rect 447692 484168 447744 484220
rect 362868 482944 362920 482996
rect 435180 482944 435232 482996
rect 506848 482944 506900 482996
rect 371148 482876 371200 482928
rect 436744 482876 436796 482928
rect 508872 482876 508924 482928
rect 513564 482876 513616 482928
rect 369216 482808 369268 482860
rect 369768 482808 369820 482860
rect 440976 482808 441028 482860
rect 512920 482808 512972 482860
rect 360844 482740 360896 482792
rect 432972 482740 433024 482792
rect 504916 482740 504968 482792
rect 323584 482400 323636 482452
rect 366916 482400 366968 482452
rect 302976 482332 303028 482384
rect 438952 482332 439004 482384
rect 198464 482264 198516 482316
rect 510896 482264 510948 482316
rect 3424 474716 3476 474768
rect 270592 474716 270644 474768
rect 227628 470568 227680 470620
rect 580172 470568 580224 470620
rect 3240 462340 3292 462392
rect 273260 462340 273312 462392
rect 445024 460164 445076 460216
rect 516416 460164 516468 460216
rect 226156 456764 226208 456816
rect 580172 456764 580224 456816
rect 373264 455404 373316 455456
rect 373908 455404 373960 455456
rect 442080 455404 442132 455456
rect 443552 455404 443604 455456
rect 3148 448536 3200 448588
rect 271880 448536 271932 448588
rect 376208 447108 376260 447160
rect 377312 447108 377364 447160
rect 442264 447108 442316 447160
rect 443460 447108 443512 447160
rect 445300 442892 445352 442944
rect 445576 442892 445628 442944
rect 467104 442892 467156 442944
rect 467748 442892 467800 442944
rect 376116 442280 376168 442332
rect 376668 442280 376720 442332
rect 377496 442280 377548 442332
rect 458824 442280 458876 442332
rect 513472 442280 513524 442332
rect 372068 442212 372120 442264
rect 460204 442212 460256 442264
rect 516600 442212 516652 442264
rect 467104 441872 467156 441924
rect 516692 441872 516744 441924
rect 457444 441804 457496 441856
rect 516968 441804 517020 441856
rect 445300 441736 445352 441788
rect 513380 441736 513432 441788
rect 445208 441668 445260 441720
rect 516508 441668 516560 441720
rect 376116 441600 376168 441652
rect 516232 441600 516284 441652
rect 516140 441532 516192 441584
rect 524420 441532 524472 441584
rect 445116 441328 445168 441380
rect 446312 441328 446364 441380
rect 446312 440376 446364 440428
rect 447876 440376 447928 440428
rect 444472 440308 444524 440360
rect 371240 440240 371292 440292
rect 371424 440240 371476 440292
rect 445576 440240 445628 440292
rect 447508 440240 447560 440292
rect 447784 440240 447836 440292
rect 513748 440240 513800 440292
rect 516876 439084 516928 439136
rect 517704 439084 517756 439136
rect 444196 439016 444248 439068
rect 447140 439016 447192 439068
rect 371792 438880 371844 438932
rect 372160 438880 372212 438932
rect 378876 438880 378928 438932
rect 516140 438880 516192 438932
rect 529940 438880 529992 438932
rect 371608 438132 371660 438184
rect 378232 438132 378284 438184
rect 444656 437928 444708 437980
rect 446036 437928 446088 437980
rect 516232 437520 516284 437572
rect 524420 437520 524472 437572
rect 378232 437452 378284 437504
rect 378968 437452 379020 437504
rect 371700 437384 371752 437436
rect 372160 437384 372212 437436
rect 371792 437316 371844 437368
rect 377036 437316 377088 437368
rect 378048 437316 378100 437368
rect 371608 437248 371660 437300
rect 380164 437452 380216 437504
rect 399484 437452 399536 437504
rect 443644 437452 443696 437504
rect 444380 437452 444432 437504
rect 446036 437452 446088 437504
rect 446680 437452 446732 437504
rect 516140 437452 516192 437504
rect 528744 437452 528796 437504
rect 516508 436840 516560 436892
rect 516876 436840 516928 436892
rect 371700 436772 371752 436824
rect 374000 436772 374052 436824
rect 379244 436772 379296 436824
rect 445116 436772 445168 436824
rect 445300 436772 445352 436824
rect 378048 436704 378100 436756
rect 387064 436704 387116 436756
rect 444380 436704 444432 436756
rect 446588 436704 446640 436756
rect 516232 436228 516284 436280
rect 523040 436228 523092 436280
rect 516508 436160 516560 436212
rect 525800 436160 525852 436212
rect 371700 436024 371752 436076
rect 379152 436092 379204 436144
rect 395344 436092 395396 436144
rect 516140 436092 516192 436144
rect 527180 436092 527232 436144
rect 371608 435956 371660 436008
rect 378784 435956 378836 436008
rect 382924 435956 382976 436008
rect 516140 434800 516192 434852
rect 521660 434800 521712 434852
rect 371700 434664 371752 434716
rect 379060 434732 379112 434784
rect 393964 434732 394016 434784
rect 516232 434732 516284 434784
rect 530032 434732 530084 434784
rect 371792 434596 371844 434648
rect 376760 434596 376812 434648
rect 380164 434596 380216 434648
rect 371608 434528 371660 434580
rect 375472 434528 375524 434580
rect 381544 434528 381596 434580
rect 444472 434392 444524 434444
rect 446128 434392 446180 434444
rect 446128 433712 446180 433764
rect 446864 433712 446916 433764
rect 516140 433440 516192 433492
rect 524512 433440 524564 433492
rect 516508 433372 516560 433424
rect 528652 433372 528704 433424
rect 516232 433304 516284 433356
rect 530124 433304 530176 433356
rect 372160 433236 372212 433288
rect 377496 433236 377548 433288
rect 444472 432896 444524 432948
rect 446220 432896 446272 432948
rect 446772 432896 446824 432948
rect 371608 432624 371660 432676
rect 376944 432760 376996 432812
rect 377404 432760 377456 432812
rect 378140 432624 378192 432676
rect 378784 432624 378836 432676
rect 371700 432556 371752 432608
rect 371424 432420 371476 432472
rect 371700 432420 371752 432472
rect 371332 432352 371384 432404
rect 371332 432148 371384 432200
rect 371608 432148 371660 432200
rect 372160 432148 372212 432200
rect 372160 432012 372212 432064
rect 372436 432012 372488 432064
rect 516508 432012 516560 432064
rect 525892 432012 525944 432064
rect 516784 431944 516836 431996
rect 528560 431944 528612 431996
rect 443092 431060 443144 431112
rect 446956 431060 447008 431112
rect 372068 429156 372120 429208
rect 372528 429156 372580 429208
rect 371608 427048 371660 427100
rect 376852 427048 376904 427100
rect 445576 426844 445628 426896
rect 447416 426844 447468 426896
rect 447968 426844 448020 426896
rect 371608 426572 371660 426624
rect 375840 426572 375892 426624
rect 376116 426572 376168 426624
rect 369124 426368 369176 426420
rect 369492 426368 369544 426420
rect 371240 426368 371292 426420
rect 375380 426368 375432 426420
rect 371608 426028 371660 426080
rect 375472 426028 375524 426080
rect 376024 426028 376076 426080
rect 516784 425688 516836 425740
rect 518164 425688 518216 425740
rect 524788 425688 524840 425740
rect 372620 425008 372672 425060
rect 372988 425008 373040 425060
rect 371056 424668 371108 424720
rect 374736 424668 374788 424720
rect 516140 424532 516192 424584
rect 517796 424532 517848 424584
rect 516140 424396 516192 424448
rect 518900 424396 518952 424448
rect 520464 424396 520516 424448
rect 516232 424328 516284 424380
rect 522028 424328 522080 424380
rect 371608 423784 371660 423836
rect 374920 423784 374972 423836
rect 371608 423648 371660 423700
rect 371976 423648 372028 423700
rect 519176 423580 519228 423632
rect 520648 423580 520700 423632
rect 371240 422560 371292 422612
rect 374644 422560 374696 422612
rect 516140 422492 516192 422544
rect 519176 422492 519228 422544
rect 516416 422424 516468 422476
rect 516140 422356 516192 422408
rect 3424 422288 3476 422340
rect 273352 422288 273404 422340
rect 516324 422288 516376 422340
rect 521936 422288 521988 422340
rect 516324 421880 516376 421932
rect 517888 421880 517940 421932
rect 371148 421608 371200 421660
rect 375012 421608 375064 421660
rect 371976 421540 372028 421592
rect 374092 421540 374144 421592
rect 374828 421540 374880 421592
rect 516324 421540 516376 421592
rect 520372 421540 520424 421592
rect 516324 421132 516376 421184
rect 520648 421132 520700 421184
rect 446496 420928 446548 420980
rect 449440 420928 449492 420980
rect 520372 420928 520424 420980
rect 521752 420928 521804 420980
rect 443828 420860 443880 420912
rect 449348 420860 449400 420912
rect 371976 420724 372028 420776
rect 374276 420724 374328 420776
rect 445576 420588 445628 420640
rect 446496 420588 446548 420640
rect 516784 420180 516836 420232
rect 518256 420180 518308 420232
rect 520280 420180 520332 420232
rect 516784 419976 516836 420028
rect 518072 419976 518124 420028
rect 518992 419976 519044 420028
rect 372436 419772 372488 419824
rect 373908 419772 373960 419824
rect 374184 419772 374236 419824
rect 516324 419772 516376 419824
rect 518900 419772 518952 419824
rect 373356 419432 373408 419484
rect 374276 419432 374328 419484
rect 444472 419432 444524 419484
rect 448704 419432 448756 419484
rect 371976 419092 372028 419144
rect 374276 419092 374328 419144
rect 516508 418548 516560 418600
rect 518992 418548 519044 418600
rect 516324 418480 516376 418532
rect 519084 418480 519136 418532
rect 372160 418140 372212 418192
rect 374460 418140 374512 418192
rect 373264 418072 373316 418124
rect 371976 417392 372028 417444
rect 377312 417392 377364 417444
rect 516324 417392 516376 417444
rect 517980 417392 518032 417444
rect 516600 417324 516652 417376
rect 517704 417324 517756 417376
rect 523132 417392 523184 417444
rect 444656 417120 444708 417172
rect 445852 417120 445904 417172
rect 446496 417120 446548 417172
rect 371976 416372 372028 416424
rect 375564 416372 375616 416424
rect 516324 415760 516376 415812
rect 520556 415760 520608 415812
rect 371976 415624 372028 415676
rect 376024 415624 376076 415676
rect 377128 415624 377180 415676
rect 516508 415420 516560 415472
rect 525984 415420 526036 415472
rect 444196 414808 444248 414860
rect 447600 414808 447652 414860
rect 371976 414740 372028 414792
rect 374552 414740 374604 414792
rect 516324 414672 516376 414724
rect 519544 414672 519596 414724
rect 522120 414672 522172 414724
rect 516324 414060 516376 414112
rect 523224 414060 523276 414112
rect 371240 413992 371292 414044
rect 516508 413992 516560 414044
rect 524604 413992 524656 414044
rect 376116 413924 376168 413976
rect 377220 413924 377272 413976
rect 445484 413652 445536 413704
rect 447324 413652 447376 413704
rect 516324 413244 516376 413296
rect 520924 413244 520976 413296
rect 524696 413244 524748 413296
rect 516784 412632 516836 412684
rect 521844 412632 521896 412684
rect 445484 412564 445536 412616
rect 447692 412564 447744 412616
rect 449256 412564 449308 412616
rect 516232 412564 516284 412616
rect 372068 412496 372120 412548
rect 372896 412496 372948 412548
rect 516324 412496 516376 412548
rect 520372 412496 520424 412548
rect 371240 412088 371292 412140
rect 375656 412088 375708 412140
rect 369124 412020 369176 412072
rect 369768 412020 369820 412072
rect 500224 412020 500276 412072
rect 516140 412020 516192 412072
rect 447692 411952 447744 412004
rect 472716 411952 472768 412004
rect 497464 411952 497516 412004
rect 516416 411952 516468 412004
rect 458824 411884 458876 411936
rect 516508 411884 516560 411936
rect 472716 411272 472768 411324
rect 513380 411272 513432 411324
rect 3148 409844 3200 409896
rect 274640 409844 274692 409896
rect 436836 409776 436888 409828
rect 508964 409776 509016 409828
rect 432880 409708 432932 409760
rect 504548 409708 504600 409760
rect 441068 409640 441120 409692
rect 513012 409640 513064 409692
rect 304264 409164 304316 409216
rect 366916 409164 366968 409216
rect 304356 409096 304408 409148
rect 438860 409096 438912 409148
rect 501604 409096 501656 409148
rect 510988 409096 511040 409148
rect 431960 408484 432012 408536
rect 432880 408484 432932 408536
rect 223396 404336 223448 404388
rect 580172 404336 580224 404388
rect 387064 398080 387116 398132
rect 450084 398080 450136 398132
rect 3424 397468 3476 397520
rect 274732 397468 274784 397520
rect 395344 395972 395396 396024
rect 395988 395972 396040 396024
rect 395988 395292 396040 395344
rect 449992 395292 450044 395344
rect 393964 394612 394016 394664
rect 394608 394612 394660 394664
rect 394608 393932 394660 393984
rect 450544 393932 450596 393984
rect 446864 389172 446916 389224
rect 447416 389172 447468 389224
rect 517888 389172 517940 389224
rect 399484 388424 399536 388476
rect 400128 388424 400180 388476
rect 448704 388424 448756 388476
rect 449164 388424 449216 388476
rect 382924 387064 382976 387116
rect 383568 387064 383620 387116
rect 441712 387064 441764 387116
rect 377404 385636 377456 385688
rect 448612 385636 448664 385688
rect 380164 384276 380216 384328
rect 448520 384276 448572 384328
rect 446772 381488 446824 381540
rect 520648 381488 520700 381540
rect 446496 380128 446548 380180
rect 523224 380128 523276 380180
rect 446496 379516 446548 379568
rect 447048 379516 447100 379568
rect 222108 378156 222160 378208
rect 580172 378156 580224 378208
rect 446680 378088 446732 378140
rect 447508 378088 447560 378140
rect 516600 377408 516652 377460
rect 522028 377408 522080 377460
rect 447508 376728 447560 376780
rect 516416 376728 516468 376780
rect 516600 376728 516652 376780
rect 447968 375980 448020 376032
rect 519084 375980 519136 376032
rect 449348 373260 449400 373312
rect 520556 373260 520608 373312
rect 378784 371832 378836 371884
rect 441620 371832 441672 371884
rect 516140 371696 516192 371748
rect 519176 371696 519228 371748
rect 3424 371220 3476 371272
rect 276020 371220 276072 371272
rect 446496 371220 446548 371272
rect 516140 371220 516192 371272
rect 506480 370472 506532 370524
rect 513380 370472 513432 370524
rect 381544 369860 381596 369912
rect 382188 369860 382240 369912
rect 444472 369860 444524 369912
rect 449900 369860 449952 369912
rect 516140 369792 516192 369844
rect 524788 369792 524840 369844
rect 372620 369656 372672 369708
rect 372896 369656 372948 369708
rect 371792 369520 371844 369572
rect 372620 369520 372672 369572
rect 370964 369316 371016 369368
rect 374736 369316 374788 369368
rect 377588 369316 377640 369368
rect 374000 369248 374052 369300
rect 441620 369248 441672 369300
rect 375288 369180 375340 369232
rect 441344 369180 441396 369232
rect 372620 369112 372672 369164
rect 442264 369112 442316 369164
rect 447876 369112 447928 369164
rect 513748 369112 513800 369164
rect 371424 368500 371476 368552
rect 375288 368500 375340 368552
rect 516140 368364 516192 368416
rect 517796 368364 517848 368416
rect 389088 367888 389140 367940
rect 441620 367888 441672 367940
rect 455328 367888 455380 367940
rect 513656 367888 513708 367940
rect 390468 367820 390520 367872
rect 441344 367820 441396 367872
rect 444564 367820 444616 367872
rect 502984 367820 503036 367872
rect 513748 367820 513800 367872
rect 370596 367752 370648 367804
rect 374644 367752 374696 367804
rect 377496 367752 377548 367804
rect 516140 367752 516192 367804
rect 520464 367752 520516 367804
rect 370320 367480 370372 367532
rect 372896 367480 372948 367532
rect 371332 367140 371384 367192
rect 374000 367140 374052 367192
rect 444288 367004 444340 367056
rect 444748 367004 444800 367056
rect 447784 366936 447836 366988
rect 454040 366936 454092 366988
rect 455328 366936 455380 366988
rect 370964 366460 371016 366512
rect 374920 366460 374972 366512
rect 377036 366460 377088 366512
rect 444656 365712 444708 365764
rect 452660 365712 452712 365764
rect 444932 365644 444984 365696
rect 448704 365644 448756 365696
rect 370964 364760 371016 364812
rect 374000 364760 374052 364812
rect 375012 364760 375064 364812
rect 444196 364352 444248 364404
rect 451280 364352 451332 364404
rect 445576 364284 445628 364336
rect 450084 364284 450136 364336
rect 445116 363808 445168 363860
rect 449992 363808 450044 363860
rect 516140 363604 516192 363656
rect 521936 363604 521988 363656
rect 369124 363536 369176 363588
rect 370320 363536 370372 363588
rect 386328 362924 386380 362976
rect 387064 362924 387116 362976
rect 445116 362856 445168 362908
rect 450176 362856 450228 362908
rect 516140 362652 516192 362704
rect 517888 362652 517940 362704
rect 370964 362448 371016 362500
rect 374092 362448 374144 362500
rect 445116 361496 445168 361548
rect 448520 361496 448572 361548
rect 516784 360816 516836 360868
rect 518256 360816 518308 360868
rect 521752 360816 521804 360868
rect 516140 360680 516192 360732
rect 520648 360680 520700 360732
rect 378048 360204 378100 360256
rect 378784 360204 378836 360256
rect 379428 360204 379480 360256
rect 380164 360204 380216 360256
rect 445116 360136 445168 360188
rect 448612 360136 448664 360188
rect 376668 359252 376720 359304
rect 377404 359252 377456 359304
rect 369768 359116 369820 359168
rect 373356 359116 373408 359168
rect 516140 359116 516192 359168
rect 518900 359116 518952 359168
rect 519176 359116 519228 359168
rect 445668 358708 445720 358760
rect 497464 358708 497516 358760
rect 516140 357892 516192 357944
rect 520280 357892 520332 357944
rect 370688 357824 370740 357876
rect 373356 357824 373408 357876
rect 369768 357756 369820 357808
rect 370136 357756 370188 357808
rect 3148 357416 3200 357468
rect 277400 357416 277452 357468
rect 445576 357348 445628 357400
rect 500224 357348 500276 357400
rect 516416 357348 516468 357400
rect 518072 357348 518124 357400
rect 445484 357280 445536 357332
rect 458824 357280 458876 357332
rect 370964 356736 371016 356788
rect 374184 356736 374236 356788
rect 516140 355580 516192 355632
rect 518992 355580 519044 355632
rect 370964 355512 371016 355564
rect 374276 355512 374328 355564
rect 445024 355308 445076 355360
rect 457444 355308 457496 355360
rect 516140 354492 516192 354544
rect 519084 354492 519136 354544
rect 370964 354424 371016 354476
rect 373264 354424 373316 354476
rect 445576 354016 445628 354068
rect 448428 354016 448480 354068
rect 449256 354016 449308 354068
rect 445116 353812 445168 353864
rect 446128 353812 446180 353864
rect 447876 353812 447928 353864
rect 446220 353336 446272 353388
rect 447968 353336 448020 353388
rect 444656 353268 444708 353320
rect 449164 353268 449216 353320
rect 445576 352588 445628 352640
rect 446036 352588 446088 352640
rect 454040 352588 454092 352640
rect 445576 352452 445628 352504
rect 447140 352452 447192 352504
rect 448612 352452 448664 352504
rect 502984 352520 503036 352572
rect 370872 352112 370924 352164
rect 374368 352112 374420 352164
rect 445576 351908 445628 351960
rect 447508 351908 447560 351960
rect 516140 351840 516192 351892
rect 523132 351840 523184 351892
rect 444380 351364 444432 351416
rect 446496 351364 446548 351416
rect 370688 351160 370740 351212
rect 377128 351160 377180 351212
rect 370596 350888 370648 350940
rect 372620 350888 372672 350940
rect 523132 350548 523184 350600
rect 524788 350548 524840 350600
rect 443828 350480 443880 350532
rect 444380 350480 444432 350532
rect 445484 350208 445536 350260
rect 447416 350208 447468 350260
rect 370964 349800 371016 349852
rect 375564 349800 375616 349852
rect 377220 349800 377272 349852
rect 516600 349800 516652 349852
rect 517704 349800 517756 349852
rect 525984 349800 526036 349852
rect 445944 349664 445996 349716
rect 446772 349664 446824 349716
rect 516140 348780 516192 348832
rect 520556 348780 520608 348832
rect 370964 348644 371016 348696
rect 376024 348644 376076 348696
rect 441896 347692 441948 347744
rect 443276 347692 443328 347744
rect 445852 347692 445904 347744
rect 446312 347692 446364 347744
rect 521016 347692 521068 347744
rect 524604 347692 524656 347744
rect 370504 347148 370556 347200
rect 375564 347148 375616 347200
rect 376116 347148 376168 347200
rect 516140 347012 516192 347064
rect 521016 347012 521068 347064
rect 444380 346672 444432 346724
rect 446404 346672 446456 346724
rect 445116 346604 445168 346656
rect 446220 346604 446272 346656
rect 516232 346332 516284 346384
rect 523224 346332 523276 346384
rect 370964 346264 371016 346316
rect 374460 346264 374512 346316
rect 516140 346264 516192 346316
rect 519544 346264 519596 346316
rect 522028 346264 522080 346316
rect 370228 345176 370280 345228
rect 373080 345176 373132 345228
rect 3332 345040 3384 345092
rect 277492 345040 277544 345092
rect 516140 344292 516192 344344
rect 519636 344292 519688 344344
rect 521844 344292 521896 344344
rect 445484 344156 445536 344208
rect 447324 344156 447376 344208
rect 370964 343952 371016 344004
rect 375656 343952 375708 344004
rect 444380 343884 444432 343936
rect 449348 343884 449400 343936
rect 514760 343544 514812 343596
rect 524696 343544 524748 343596
rect 370964 342864 371016 342916
rect 372712 342864 372764 342916
rect 377312 342864 377364 342916
rect 443644 342252 443696 342304
rect 444656 342252 444708 342304
rect 445116 342252 445168 342304
rect 447048 342252 447100 342304
rect 447600 342184 447652 342236
rect 514760 342048 514812 342100
rect 516140 341708 516192 341760
rect 520372 341708 520424 341760
rect 441620 340892 441672 340944
rect 447600 340892 447652 340944
rect 446404 340824 446456 340876
rect 516416 340824 516468 340876
rect 472624 340756 472676 340808
rect 513380 340756 513432 340808
rect 445484 340552 445536 340604
rect 447232 340552 447284 340604
rect 444564 339464 444616 339516
rect 471244 339464 471296 339516
rect 472624 339464 472676 339516
rect 368940 339192 368992 339244
rect 369308 339192 369360 339244
rect 506848 338036 506900 338088
rect 507768 338036 507820 338088
rect 513472 338036 513524 338088
rect 512920 337696 512972 337748
rect 514760 337696 514812 337748
rect 322204 337424 322256 337476
rect 366916 337424 366968 337476
rect 431224 337424 431276 337476
rect 438952 337424 439004 337476
rect 300768 337356 300820 337408
rect 510896 337356 510948 337408
rect 246948 330488 247000 330540
rect 331220 330488 331272 330540
rect 41328 327700 41380 327752
rect 258080 327700 258132 327752
rect 443644 326272 443696 326324
rect 444196 326272 444248 326324
rect 523040 326340 523092 326392
rect 219348 324300 219400 324352
rect 579620 324300 579672 324352
rect 378048 322192 378100 322244
rect 525892 322192 525944 322244
rect 377404 321580 377456 321632
rect 378048 321580 378100 321632
rect 373356 318860 373408 318912
rect 373816 318860 373868 318912
rect 3424 318792 3476 318844
rect 278780 318792 278832 318844
rect 441988 318792 442040 318844
rect 443276 318792 443328 318844
rect 395344 318724 395396 318776
rect 395988 318724 396040 318776
rect 395344 318044 395396 318096
rect 521660 318044 521712 318096
rect 379428 315256 379480 315308
rect 524512 315256 524564 315308
rect 378784 314644 378836 314696
rect 379428 314644 379480 314696
rect 373264 313896 373316 313948
rect 446220 313896 446272 313948
rect 220636 311856 220688 311908
rect 580172 311856 580224 311908
rect 385776 310088 385828 310140
rect 386328 310088 386380 310140
rect 386328 309748 386380 309800
rect 527180 309748 527232 309800
rect 376024 309068 376076 309120
rect 441896 309068 441948 309120
rect 444564 309068 444616 309120
rect 244464 307164 244516 307216
rect 396724 307164 396776 307216
rect 241888 307096 241940 307148
rect 461584 307096 461636 307148
rect 239312 307028 239364 307080
rect 526444 307028 526496 307080
rect 248696 306008 248748 306060
rect 295984 306008 296036 306060
rect 171048 305940 171100 305992
rect 253756 305940 253808 305992
rect 246120 305872 246172 305924
rect 359464 305872 359516 305924
rect 106188 305804 106240 305856
rect 256240 305804 256292 305856
rect 243544 305736 243596 305788
rect 429200 305736 429252 305788
rect 228272 305668 228324 305720
rect 582380 305668 582432 305720
rect 226616 305600 226668 305652
rect 582472 305600 582524 305652
rect 3240 304988 3292 305040
rect 280896 304988 280948 305040
rect 233148 304784 233200 304836
rect 251180 304784 251232 304836
rect 241060 304716 241112 304768
rect 494060 304716 494112 304768
rect 238484 304648 238536 304700
rect 558920 304648 558972 304700
rect 232596 304580 232648 304632
rect 580264 304580 580316 304632
rect 230848 304512 230900 304564
rect 580356 304512 580408 304564
rect 224960 304444 225012 304496
rect 580540 304444 580592 304496
rect 224040 304376 224092 304428
rect 580448 304376 580500 304428
rect 222384 304308 222436 304360
rect 580632 304308 580684 304360
rect 220728 304240 220780 304292
rect 580724 304240 580776 304292
rect 262220 303220 262272 303272
rect 262772 303220 262824 303272
rect 274640 303220 274692 303272
rect 275468 303220 275520 303272
rect 277400 303220 277452 303272
rect 278044 303220 278096 303272
rect 212172 303152 212224 303204
rect 536104 303152 536156 303204
rect 207112 303084 207164 303136
rect 533344 303084 533396 303136
rect 204628 303016 204680 303068
rect 530584 303016 530636 303068
rect 43444 302948 43496 303000
rect 296076 302948 296128 303000
rect 28264 302880 28316 302932
rect 285956 302880 286008 302932
rect 29644 302812 29696 302864
rect 288532 302812 288584 302864
rect 299480 302812 299532 302864
rect 300768 302812 300820 302864
rect 32404 302744 32456 302796
rect 293592 302744 293644 302796
rect 26884 302676 26936 302728
rect 295248 302676 295300 302728
rect 4804 302608 4856 302660
rect 291016 302608 291068 302660
rect 211344 302540 211396 302592
rect 522304 302540 522356 302592
rect 208860 302472 208912 302524
rect 520924 302472 520976 302524
rect 202052 302404 202104 302456
rect 525064 302404 525116 302456
rect 296996 302336 297048 302388
rect 297824 302268 297876 302320
rect 298652 302200 298704 302252
rect 305644 302200 305696 302252
rect 307024 302268 307076 302320
rect 309784 302200 309836 302252
rect 229192 302064 229244 302116
rect 230388 302064 230440 302116
rect 199384 301588 199436 301640
rect 284208 301588 284260 301640
rect 210516 301520 210568 301572
rect 301504 301520 301556 301572
rect 215576 301452 215628 301504
rect 312544 301452 312596 301504
rect 206284 301384 206336 301436
rect 318064 301384 318116 301436
rect 201224 301316 201276 301368
rect 313924 301316 313976 301368
rect 152464 301248 152516 301300
rect 287612 301248 287664 301300
rect 156604 301180 156656 301232
rect 294420 301180 294472 301232
rect 148324 301112 148376 301164
rect 292764 301112 292816 301164
rect 10324 301044 10376 301096
rect 281724 301044 281776 301096
rect 214748 300976 214800 301028
rect 519544 300976 519596 301028
rect 202880 300908 202932 300960
rect 582472 300908 582524 300960
rect 200396 300840 200448 300892
rect 582380 300840 582432 300892
rect 219808 300228 219860 300280
rect 220636 300228 220688 300280
rect 233424 300228 233476 300280
rect 234436 300228 234488 300280
rect 237656 300228 237708 300280
rect 238576 300228 238628 300280
rect 240140 300228 240192 300280
rect 241336 300228 241388 300280
rect 205456 300160 205508 300212
rect 311164 300160 311216 300212
rect 203708 300092 203760 300144
rect 316684 300092 316736 300144
rect 155224 300024 155276 300076
rect 284852 300024 284904 300076
rect 159364 299956 159416 300008
rect 289084 299956 289136 300008
rect 157984 299888 158036 299940
rect 291476 299888 291528 299940
rect 151084 299820 151136 299872
rect 289820 299820 289872 299872
rect 371424 299820 371476 299872
rect 375288 299820 375340 299872
rect 11704 299752 11756 299804
rect 286508 299752 286560 299804
rect 213368 299684 213420 299736
rect 515404 299684 515456 299736
rect 210056 299616 210108 299668
rect 518164 299616 518216 299668
rect 208216 299548 208268 299600
rect 526444 299548 526496 299600
rect 218520 299480 218572 299532
rect 580172 299480 580224 299532
rect 214012 299412 214064 299464
rect 198464 298528 198516 298580
rect 3884 298460 3936 298512
rect 214012 299276 214064 299328
rect 214564 299276 214616 299328
rect 214656 299276 214708 299328
rect 216036 299276 216088 299328
rect 216864 299276 216916 299328
rect 216956 299276 217008 299328
rect 217600 299276 217652 299328
rect 3424 298392 3476 298444
rect 3516 298324 3568 298376
rect 224408 299276 224460 299328
rect 282644 299412 282696 299464
rect 283472 299412 283524 299464
rect 279700 299276 279752 299328
rect 282276 299276 282328 299328
rect 282644 299276 282696 299328
rect 283012 299276 283064 299328
rect 283472 299276 283524 299328
rect 375932 299072 375984 299124
rect 376668 299072 376720 299124
rect 382280 298800 382332 298852
rect 394608 298800 394660 298852
rect 516784 298800 516836 298852
rect 379428 298732 379480 298784
rect 383568 298732 383620 298784
rect 516600 298732 516652 298784
rect 429844 298528 429896 298580
rect 507768 298460 507820 298512
rect 514208 298460 514260 298512
rect 382188 298392 382240 298444
rect 516692 298392 516744 298444
rect 375932 298324 375984 298376
rect 516508 298324 516560 298376
rect 580356 298256 580408 298308
rect 580448 298188 580500 298240
rect 580264 298120 580316 298172
rect 441896 298052 441948 298104
rect 442448 298052 442500 298104
rect 445300 298052 445352 298104
rect 445668 298052 445720 298104
rect 371332 297984 371384 298036
rect 375196 297984 375248 298036
rect 445116 297984 445168 298036
rect 445576 297984 445628 298036
rect 507860 297848 507912 297900
rect 513748 297848 513800 297900
rect 442448 297576 442500 297628
rect 444380 297508 444432 297560
rect 446128 297508 446180 297560
rect 303068 297440 303120 297492
rect 369400 297440 369452 297492
rect 443276 297440 443328 297492
rect 444288 297440 444340 297492
rect 516324 297508 516376 297560
rect 302884 297372 302936 297424
rect 369860 297372 369912 297424
rect 375196 297372 375248 297424
rect 513380 297372 513432 297424
rect 448428 297304 448480 297356
rect 517152 297304 517204 297356
rect 445392 297236 445444 297288
rect 514116 297236 514168 297288
rect 445116 297168 445168 297220
rect 513288 297168 513340 297220
rect 444932 297100 444984 297152
rect 513932 297100 513984 297152
rect 444748 297032 444800 297084
rect 513840 297032 513892 297084
rect 445668 296964 445720 297016
rect 516416 296964 516468 297016
rect 444288 296896 444340 296948
rect 516232 296896 516284 296948
rect 442264 296828 442316 296880
rect 516140 296828 516192 296880
rect 371792 296760 371844 296812
rect 425704 296760 425756 296812
rect 441712 296760 441764 296812
rect 375104 296692 375156 296744
rect 513380 296692 513432 296744
rect 371240 296624 371292 296676
rect 389088 296624 389140 296676
rect 390468 296556 390520 296608
rect 513380 296556 513432 296608
rect 517244 296556 517296 296608
rect 378876 296488 378928 296540
rect 443276 296488 443328 296540
rect 444380 296488 444432 296540
rect 446036 296488 446088 296540
rect 389088 296420 389140 296472
rect 513472 296420 513524 296472
rect 347688 296148 347740 296200
rect 369400 296148 369452 296200
rect 371240 296148 371292 296200
rect 375288 296148 375340 296200
rect 391940 296148 391992 296200
rect 372344 296080 372396 296132
rect 390468 296080 390520 296132
rect 400680 296080 400732 296132
rect 443644 296080 443696 296132
rect 358084 296012 358136 296064
rect 371424 296012 371476 296064
rect 388444 296012 388496 296064
rect 441896 296012 441948 296064
rect 372160 295944 372212 295996
rect 442080 295944 442132 295996
rect 445208 295944 445260 295996
rect 428464 295876 428516 295928
rect 441712 295876 441764 295928
rect 517244 295944 517296 295996
rect 528836 295944 528888 295996
rect 359464 295808 359516 295860
rect 369860 295808 369912 295860
rect 391940 295808 391992 295860
rect 393228 295808 393280 295860
rect 513564 295808 513616 295860
rect 513656 295468 513708 295520
rect 379244 295400 379296 295452
rect 400680 295400 400732 295452
rect 302792 295332 302844 295384
rect 320824 295332 320876 295384
rect 378968 295332 379020 295384
rect 388444 295332 388496 295384
rect 371332 295264 371384 295316
rect 378876 295264 378928 295316
rect 516140 295264 516192 295316
rect 529940 295264 529992 295316
rect 371700 295196 371752 295248
rect 378968 295196 379020 295248
rect 445392 295196 445444 295248
rect 448612 295196 448664 295248
rect 516324 295196 516376 295248
rect 528744 295196 528796 295248
rect 445484 295128 445536 295180
rect 447508 295128 447560 295180
rect 516232 295128 516284 295180
rect 524420 295128 524472 295180
rect 447508 294584 447560 294636
rect 456064 294584 456116 294636
rect 448612 293972 448664 294024
rect 449256 293972 449308 294024
rect 371240 293904 371292 293956
rect 400128 293904 400180 293956
rect 516232 293904 516284 293956
rect 525800 293904 525852 293956
rect 371332 293836 371384 293888
rect 379244 293836 379296 293888
rect 516140 293836 516192 293888
rect 523040 293836 523092 293888
rect 371240 292476 371292 292528
rect 385776 292476 385828 292528
rect 516324 292476 516376 292528
rect 516600 292476 516652 292528
rect 530032 292476 530084 292528
rect 516140 292408 516192 292460
rect 527180 292408 527232 292460
rect 516232 292340 516284 292392
rect 521660 292340 521712 292392
rect 513748 291864 513800 291916
rect 514024 291864 514076 291916
rect 371700 291796 371752 291848
rect 378232 291796 378284 291848
rect 379428 291796 379480 291848
rect 386328 291796 386380 291848
rect 395344 291796 395396 291848
rect 372252 291728 372304 291780
rect 372436 291728 372488 291780
rect 371700 291184 371752 291236
rect 385684 291184 385736 291236
rect 386328 291184 386380 291236
rect 380900 291116 380952 291168
rect 382188 291116 382240 291168
rect 516324 291116 516376 291168
rect 516784 291116 516836 291168
rect 530124 291116 530176 291168
rect 516232 291048 516284 291100
rect 516692 291048 516744 291100
rect 528652 291048 528704 291100
rect 371332 290640 371384 290692
rect 371884 290640 371936 290692
rect 371700 290504 371752 290556
rect 380900 290504 380952 290556
rect 371792 290436 371844 290488
rect 382280 290436 382332 290488
rect 445484 290368 445536 290420
rect 447416 290368 447468 290420
rect 447968 290368 448020 290420
rect 170404 289824 170456 289876
rect 197360 289824 197412 289876
rect 444288 289824 444340 289876
rect 447876 289824 447928 289876
rect 376024 289756 376076 289808
rect 377404 289756 377456 289808
rect 378140 289756 378192 289808
rect 378784 289756 378836 289808
rect 516324 289756 516376 289808
rect 516508 289756 516560 289808
rect 528560 289756 528612 289808
rect 516232 289688 516284 289740
rect 525892 289688 525944 289740
rect 516140 289620 516192 289672
rect 524512 289620 524564 289672
rect 302240 289212 302292 289264
rect 304356 289212 304408 289264
rect 371700 289212 371752 289264
rect 376024 289212 376076 289264
rect 371240 289076 371292 289128
rect 378140 289076 378192 289128
rect 371700 288532 371752 288584
rect 375932 288532 375984 288584
rect 445944 287444 445996 287496
rect 446680 287444 446732 287496
rect 443184 287104 443236 287156
rect 447784 287104 447836 287156
rect 178684 287036 178736 287088
rect 198556 287036 198608 287088
rect 302240 286492 302292 286544
rect 304264 286492 304316 286544
rect 371148 286356 371200 286408
rect 371608 286356 371660 286408
rect 371516 286288 371568 286340
rect 377404 286288 377456 286340
rect 371976 285676 372028 285728
rect 374552 285676 374604 285728
rect 444748 284792 444800 284844
rect 446404 284792 446456 284844
rect 372252 284316 372304 284368
rect 375380 284316 375432 284368
rect 369216 283568 369268 283620
rect 369676 283568 369728 283620
rect 371516 283568 371568 283620
rect 376760 283568 376812 283620
rect 376944 283568 376996 283620
rect 369124 283296 369176 283348
rect 369400 283296 369452 283348
rect 174544 282888 174596 282940
rect 197360 282888 197412 282940
rect 302792 282888 302844 282940
rect 353944 282888 353996 282940
rect 445852 282888 445904 282940
rect 446588 282888 446640 282940
rect 377588 282820 377640 282872
rect 378048 282820 378100 282872
rect 425704 282820 425756 282872
rect 444380 282820 444432 282872
rect 446220 282820 446272 282872
rect 371700 282276 371752 282328
rect 375472 282276 375524 282328
rect 377680 282276 377732 282328
rect 371608 282208 371660 282260
rect 375840 282208 375892 282260
rect 376852 282208 376904 282260
rect 371516 282140 371568 282192
rect 378048 282140 378100 282192
rect 160100 281528 160152 281580
rect 197912 281528 197964 281580
rect 516140 281528 516192 281580
rect 524512 281528 524564 281580
rect 377496 281460 377548 281512
rect 378048 281460 378100 281512
rect 428464 281460 428516 281512
rect 444748 281256 444800 281308
rect 445760 281256 445812 281308
rect 446772 281256 446824 281308
rect 369216 280848 369268 280900
rect 369400 280848 369452 280900
rect 371516 280780 371568 280832
rect 378048 280780 378100 280832
rect 445484 280576 445536 280628
rect 447324 280576 447376 280628
rect 448060 280576 448112 280628
rect 516140 280440 516192 280492
rect 518900 280440 518952 280492
rect 516232 280168 516284 280220
rect 521660 280168 521712 280220
rect 371424 279420 371476 279472
rect 377036 279420 377088 279472
rect 517796 279420 517848 279472
rect 521936 279420 521988 279472
rect 371608 279352 371660 279404
rect 374000 279352 374052 279404
rect 374736 279352 374788 279404
rect 516140 278808 516192 278860
rect 523132 278808 523184 278860
rect 175924 278740 175976 278792
rect 197544 278740 197596 278792
rect 302424 278740 302476 278792
rect 356704 278740 356756 278792
rect 516232 278740 516284 278792
rect 524420 278740 524472 278792
rect 376116 278672 376168 278724
rect 377036 278672 377088 278724
rect 516140 278672 516192 278724
rect 516416 278672 516468 278724
rect 371608 278264 371660 278316
rect 374092 278264 374144 278316
rect 374828 278264 374880 278316
rect 516692 277856 516744 277908
rect 518256 277856 518308 277908
rect 518256 277448 518308 277500
rect 519268 277448 519320 277500
rect 181444 277380 181496 277432
rect 197360 277380 197412 277432
rect 516416 277380 516468 277432
rect 521752 277380 521804 277432
rect 516140 276904 516192 276956
rect 516416 276904 516468 276956
rect 516140 276768 516192 276820
rect 519176 276768 519228 276820
rect 516692 276292 516744 276344
rect 518072 276292 518124 276344
rect 520280 276292 520332 276344
rect 372436 276224 372488 276276
rect 373908 276224 373960 276276
rect 371424 276156 371476 276208
rect 374644 276156 374696 276208
rect 519176 276088 519228 276140
rect 520464 276088 520516 276140
rect 302792 276020 302844 276072
rect 358176 276020 358228 276072
rect 516324 276020 516376 276072
rect 521936 276020 521988 276072
rect 371608 275748 371660 275800
rect 374184 275748 374236 275800
rect 372804 275340 372856 275392
rect 373264 275340 373316 275392
rect 372160 275204 372212 275256
rect 373264 275204 373316 275256
rect 374276 275204 374328 275256
rect 516140 275204 516192 275256
rect 519084 275204 519136 275256
rect 516324 275136 516376 275188
rect 520556 275136 520608 275188
rect 188344 274660 188396 274712
rect 197544 274660 197596 274712
rect 516140 274660 516192 274712
rect 518348 274660 518400 274712
rect 373356 274592 373408 274644
rect 374184 274592 374236 274644
rect 516692 274048 516744 274100
rect 517612 274048 517664 274100
rect 519176 274048 519228 274100
rect 371608 273572 371660 273624
rect 374000 273572 374052 273624
rect 374368 273572 374420 273624
rect 180064 273232 180116 273284
rect 197360 273232 197412 273284
rect 302700 273232 302752 273284
rect 360568 273232 360620 273284
rect 371516 273232 371568 273284
rect 372620 273232 372672 273284
rect 372896 273232 372948 273284
rect 517520 273232 517572 273284
rect 518256 273232 518308 273284
rect 444564 273164 444616 273216
rect 447140 273164 447192 273216
rect 516140 273164 516192 273216
rect 524788 273164 524840 273216
rect 528652 273164 528704 273216
rect 516324 272484 516376 272536
rect 517888 272484 517940 272536
rect 516140 271872 516192 271924
rect 525892 271872 525944 271924
rect 371884 271804 371936 271856
rect 372252 271804 372304 271856
rect 377220 271804 377272 271856
rect 371700 271736 371752 271788
rect 377128 271736 377180 271788
rect 371792 271668 371844 271720
rect 372160 271668 372212 271720
rect 376208 271668 376260 271720
rect 516140 271192 516192 271244
rect 521016 271192 521068 271244
rect 524604 271192 524656 271244
rect 516324 271124 516376 271176
rect 521844 271124 521896 271176
rect 522028 271124 522080 271176
rect 372528 270580 372580 270632
rect 375564 270580 375616 270632
rect 186964 270512 187016 270564
rect 197544 270512 197596 270564
rect 371792 270444 371844 270496
rect 372068 270444 372120 270496
rect 374460 270444 374512 270496
rect 516140 270172 516192 270224
rect 519636 270172 519688 270224
rect 523040 270172 523092 270224
rect 371424 269764 371476 269816
rect 377312 270036 377364 270088
rect 441620 270036 441672 270088
rect 445484 269764 445536 269816
rect 447232 269764 447284 269816
rect 516324 269492 516376 269544
rect 520648 269492 520700 269544
rect 193864 269288 193916 269340
rect 198464 269288 198516 269340
rect 516140 269084 516192 269136
rect 525800 269084 525852 269136
rect 371884 269016 371936 269068
rect 375656 269016 375708 269068
rect 471060 269016 471112 269068
rect 471244 269016 471296 269068
rect 513380 269016 513432 269068
rect 371976 268948 372028 269000
rect 373080 268948 373132 269000
rect 513288 268948 513340 269000
rect 514760 268948 514812 269000
rect 516140 268608 516192 268660
rect 520372 268608 520424 268660
rect 486424 268540 486476 268592
rect 516508 268540 516560 268592
rect 445484 268472 445536 268524
rect 445760 268472 445812 268524
rect 471060 268472 471112 268524
rect 476764 268472 476816 268524
rect 516416 268472 516468 268524
rect 303344 268404 303396 268456
rect 369952 268404 370004 268456
rect 457444 268404 457496 268456
rect 516600 268404 516652 268456
rect 303252 268336 303304 268388
rect 370688 268336 370740 268388
rect 444564 268336 444616 268388
rect 445484 268336 445536 268388
rect 449348 268336 449400 268388
rect 516784 268336 516836 268388
rect 369952 268268 370004 268320
rect 370228 268268 370280 268320
rect 369124 268200 369176 268252
rect 369032 267996 369084 268048
rect 2964 267656 3016 267708
rect 10324 267656 10376 267708
rect 449164 267656 449216 267708
rect 516232 267656 516284 267708
rect 303160 266976 303212 267028
rect 370596 266976 370648 267028
rect 184204 266364 184256 266416
rect 197636 266364 197688 266416
rect 362868 266296 362920 266348
rect 431776 266296 431828 266348
rect 434904 266296 434956 266348
rect 364892 266228 364944 266280
rect 431868 266228 431920 266280
rect 436928 266228 436980 266280
rect 503720 266296 503772 266348
rect 504916 266296 504968 266348
rect 506848 266296 506900 266348
rect 507768 266296 507820 266348
rect 513748 266296 513800 266348
rect 353944 266160 353996 266212
rect 368940 266160 368992 266212
rect 369124 266160 369176 266212
rect 370228 266160 370280 266212
rect 429844 266160 429896 266212
rect 438860 266160 438912 266212
rect 508872 266228 508924 266280
rect 509148 266228 509200 266280
rect 513472 266228 513524 266280
rect 307024 266092 307076 266144
rect 366916 266092 366968 266144
rect 360200 265684 360252 265736
rect 360936 265684 360988 265736
rect 431960 265684 432012 265736
rect 432880 265684 432932 265736
rect 503720 265684 503772 265736
rect 370228 265616 370280 265668
rect 440608 265616 440660 265668
rect 441068 265616 441120 265668
rect 512644 265616 512696 265668
rect 182824 264936 182876 264988
rect 197360 264936 197412 264988
rect 502984 264936 503036 264988
rect 510896 264936 510948 264988
rect 302700 264868 302752 264920
rect 358084 264868 358136 264920
rect 302884 264188 302936 264240
rect 369492 264188 369544 264240
rect 181536 262216 181588 262268
rect 197360 262216 197412 262268
rect 302332 262148 302384 262200
rect 359464 262148 359516 262200
rect 180156 260856 180208 260908
rect 197360 260856 197412 260908
rect 357348 260108 357400 260160
rect 370504 260108 370556 260160
rect 313188 258680 313240 258732
rect 347688 258680 347740 258732
rect 442080 258680 442132 258732
rect 178776 258068 178828 258120
rect 197360 258068 197412 258120
rect 302608 258068 302660 258120
rect 313188 258068 313240 258120
rect 196624 256708 196676 256760
rect 198372 256708 198424 256760
rect 302792 255960 302844 256012
rect 357348 255960 357400 256012
rect 357348 255280 357400 255332
rect 441712 255280 441764 255332
rect 195244 253920 195296 253972
rect 198004 253920 198056 253972
rect 192576 251200 192628 251252
rect 197912 251200 197964 251252
rect 302976 251200 303028 251252
rect 307668 251200 307720 251252
rect 441804 251200 441856 251252
rect 303344 250452 303396 250504
rect 370412 250452 370464 250504
rect 191196 249772 191248 249824
rect 198096 249772 198148 249824
rect 370412 249024 370464 249076
rect 388444 249024 388496 249076
rect 441896 249024 441948 249076
rect 302792 248412 302844 248464
rect 370412 248412 370464 248464
rect 444380 247868 444432 247920
rect 445208 247868 445260 247920
rect 371056 247664 371108 247716
rect 444380 247664 444432 247716
rect 446680 247664 446732 247716
rect 521936 247664 521988 247716
rect 177396 247052 177448 247104
rect 197544 247052 197596 247104
rect 370504 247052 370556 247104
rect 371056 247052 371108 247104
rect 340328 246304 340380 246356
rect 400864 246304 400916 246356
rect 441988 246304 442040 246356
rect 302516 245624 302568 245676
rect 340328 245624 340380 245676
rect 340788 245624 340840 245676
rect 312544 245556 312596 245608
rect 580172 245556 580224 245608
rect 446496 243516 446548 243568
rect 446864 243516 446916 243568
rect 517796 243516 517848 243568
rect 517980 243516 518032 243568
rect 171784 242904 171836 242956
rect 197544 242904 197596 242956
rect 303252 242904 303304 242956
rect 443552 242904 443604 242956
rect 377404 242836 377456 242888
rect 377772 242836 377824 242888
rect 444472 242836 444524 242888
rect 444932 242836 444984 242888
rect 342904 242156 342956 242208
rect 377772 242156 377824 242208
rect 195336 241476 195388 241528
rect 198280 241476 198332 241528
rect 444564 241408 444616 241460
rect 444840 241408 444892 241460
rect 446496 241408 446548 241460
rect 446772 241408 446824 241460
rect 304264 240728 304316 240780
rect 374552 240728 374604 240780
rect 406384 240728 406436 240780
rect 446496 240728 446548 240780
rect 519176 240728 519228 240780
rect 406384 240116 406436 240168
rect 444564 240116 444616 240168
rect 444656 240048 444708 240100
rect 445208 240048 445260 240100
rect 445208 239368 445260 239420
rect 517888 239368 517940 239420
rect 171876 238756 171928 238808
rect 197544 238756 197596 238808
rect 443644 238348 443696 238400
rect 444288 238348 444340 238400
rect 444288 238008 444340 238060
rect 523132 238008 523184 238060
rect 196716 237736 196768 237788
rect 198464 237736 198516 237788
rect 378232 236648 378284 236700
rect 443184 236648 443236 236700
rect 446588 236648 446640 236700
rect 519084 236648 519136 236700
rect 302792 235968 302844 236020
rect 375472 235968 375524 236020
rect 378232 235968 378284 236020
rect 447968 235220 448020 235272
rect 521752 235220 521804 235272
rect 522028 235220 522080 235272
rect 171968 234608 172020 234660
rect 197544 234608 197596 234660
rect 516232 234540 516284 234592
rect 518900 234540 518952 234592
rect 376668 233860 376720 233912
rect 385684 233860 385736 233912
rect 443276 233860 443328 233912
rect 445300 233860 445352 233912
rect 528652 233860 528704 233912
rect 172060 233248 172112 233300
rect 197360 233248 197412 233300
rect 302700 233248 302752 233300
rect 375564 233248 375616 233300
rect 376668 233248 376720 233300
rect 449256 233248 449308 233300
rect 516232 233248 516284 233300
rect 516600 233248 516652 233300
rect 447876 233180 447928 233232
rect 448152 233180 448204 233232
rect 516416 233180 516468 233232
rect 519268 233180 519320 233232
rect 448152 231820 448204 231872
rect 516416 231820 516468 231872
rect 375656 231072 375708 231124
rect 380900 231072 380952 231124
rect 443368 231072 443420 231124
rect 444932 231072 444984 231124
rect 521844 231072 521896 231124
rect 302792 230460 302844 230512
rect 375656 230460 375708 230512
rect 444840 230392 444892 230444
rect 445116 230392 445168 230444
rect 371148 229712 371200 229764
rect 444840 229712 444892 229764
rect 446404 229712 446456 229764
rect 520556 229712 520608 229764
rect 174636 229100 174688 229152
rect 197360 229100 197412 229152
rect 517704 228692 517756 228744
rect 518256 228692 518308 228744
rect 448060 228420 448112 228472
rect 517704 228420 517756 228472
rect 445392 228352 445444 228404
rect 524604 228352 524656 228404
rect 441804 228284 441856 228336
rect 442356 228284 442408 228336
rect 447876 227740 447928 227792
rect 448060 227740 448112 227792
rect 302792 227672 302844 227724
rect 382280 227672 382332 227724
rect 382280 226992 382332 227044
rect 394148 226992 394200 227044
rect 516232 226788 516284 226840
rect 520464 226788 520516 226840
rect 176016 226312 176068 226364
rect 197544 226312 197596 226364
rect 394148 226312 394200 226364
rect 394608 226312 394660 226364
rect 443460 226312 443512 226364
rect 447784 226312 447836 226364
rect 516232 226312 516284 226364
rect 516508 226312 516560 226364
rect 375196 226244 375248 226296
rect 441620 226244 441672 226296
rect 516140 226244 516192 226296
rect 524512 226244 524564 226296
rect 375104 226176 375156 226228
rect 441620 226108 441672 226160
rect 304908 225632 304960 225684
rect 367836 225632 367888 225684
rect 509148 225632 509200 225684
rect 514852 225632 514904 225684
rect 302976 225564 303028 225616
rect 371148 225564 371200 225616
rect 507768 225564 507820 225616
rect 512644 225564 512696 225616
rect 514944 225564 514996 225616
rect 514760 225496 514812 225548
rect 441988 225156 442040 225208
rect 442264 225156 442316 225208
rect 441896 225088 441948 225140
rect 442172 225088 442224 225140
rect 351920 225020 351972 225072
rect 375840 225020 375892 225072
rect 445944 225020 445996 225072
rect 464344 225020 464396 225072
rect 513748 225020 513800 225072
rect 177304 224952 177356 225004
rect 197360 224952 197412 225004
rect 345664 224952 345716 225004
rect 375748 224952 375800 225004
rect 445852 224952 445904 225004
rect 456064 224952 456116 225004
rect 513380 224952 513432 225004
rect 390468 224884 390520 224936
rect 441712 224884 441764 224936
rect 516140 224884 516192 224936
rect 521660 224884 521712 224936
rect 393228 224816 393280 224868
rect 441620 224816 441672 224868
rect 302884 224340 302936 224392
rect 340880 224340 340932 224392
rect 358084 224272 358136 224324
rect 369400 224272 369452 224324
rect 371332 224272 371384 224324
rect 444472 224272 444524 224324
rect 445576 224272 445628 224324
rect 302884 224204 302936 224256
rect 370504 224204 370556 224256
rect 378140 224204 378192 224256
rect 443184 224204 443236 224256
rect 445116 224204 445168 224256
rect 445668 224204 445720 224256
rect 302332 223932 302384 223984
rect 375932 223932 375984 223984
rect 378140 223932 378192 223984
rect 340880 223864 340932 223916
rect 342168 223864 342220 223916
rect 441804 223864 441856 223916
rect 461584 223864 461636 223916
rect 513748 223864 513800 223916
rect 170496 222844 170548 222896
rect 198188 222844 198240 222896
rect 444748 222300 444800 222352
rect 483664 222300 483716 222352
rect 445576 222232 445628 222284
rect 489184 222232 489236 222284
rect 445668 222164 445720 222216
rect 485044 222164 485096 222216
rect 302332 222096 302384 222148
rect 351920 222096 351972 222148
rect 454684 222096 454736 222148
rect 456064 222096 456116 222148
rect 516140 222096 516192 222148
rect 524420 222096 524472 222148
rect 191104 220872 191156 220924
rect 197360 220872 197412 220924
rect 370320 220872 370372 220924
rect 376024 220872 376076 220924
rect 444748 220872 444800 220924
rect 482284 220872 482336 220924
rect 445576 220804 445628 220856
rect 490564 220804 490616 220856
rect 371516 220736 371568 220788
rect 372436 220736 372488 220788
rect 376116 220736 376168 220788
rect 516140 220736 516192 220788
rect 523132 220736 523184 220788
rect 516140 219920 516192 219972
rect 517980 219920 518032 219972
rect 445668 219580 445720 219632
rect 479524 219580 479576 219632
rect 443276 219512 443328 219564
rect 444748 219512 444800 219564
rect 493324 219512 493376 219564
rect 302424 219376 302476 219428
rect 345664 219376 345716 219428
rect 445576 219444 445628 219496
rect 494704 219444 494756 219496
rect 443644 219376 443696 219428
rect 519544 219376 519596 219428
rect 580172 219376 580224 219428
rect 516140 219308 516192 219360
rect 522028 219308 522080 219360
rect 370320 218424 370372 218476
rect 374184 218424 374236 218476
rect 374828 218424 374880 218476
rect 443644 218084 443696 218136
rect 475384 218084 475436 218136
rect 192484 218016 192536 218068
rect 197544 218016 197596 218068
rect 443368 218016 443420 218068
rect 497464 218016 497516 218068
rect 370964 217336 371016 217388
rect 372988 217336 373040 217388
rect 517060 217336 517112 217388
rect 518900 217336 518952 217388
rect 445944 217268 445996 217320
rect 471244 217268 471296 217320
rect 188436 216656 188488 216708
rect 197360 216656 197412 216708
rect 372988 216656 373040 216708
rect 373540 216656 373592 216708
rect 443276 216656 443328 216708
rect 472624 216656 472676 216708
rect 516140 216588 516192 216640
rect 521936 216588 521988 216640
rect 370964 216180 371016 216232
rect 374644 216180 374696 216232
rect 303068 215908 303120 215960
rect 303528 215908 303580 215960
rect 352564 215908 352616 215960
rect 445852 215908 445904 215960
rect 468484 215908 468536 215960
rect 444472 215840 444524 215892
rect 446036 215840 446088 215892
rect 3332 215228 3384 215280
rect 199384 215228 199436 215280
rect 370688 215024 370740 215076
rect 374368 215024 374420 215076
rect 187056 213936 187108 213988
rect 197360 213936 197412 213988
rect 372804 213868 372856 213920
rect 373356 213868 373408 213920
rect 516232 213868 516284 213920
rect 518072 213868 518124 213920
rect 370964 213800 371016 213852
rect 374276 213800 374328 213852
rect 516140 213800 516192 213852
rect 520556 213800 520608 213852
rect 445116 212848 445168 212900
rect 445944 212848 445996 212900
rect 444748 212440 444800 212492
rect 486424 212440 486476 212492
rect 442724 212372 442776 212424
rect 445024 212372 445076 212424
rect 476764 212372 476816 212424
rect 445116 212304 445168 212356
rect 457444 212304 457496 212356
rect 516140 211896 516192 211948
rect 519084 211896 519136 211948
rect 370964 211556 371016 211608
rect 373448 211556 373500 211608
rect 184296 211148 184348 211200
rect 197360 211148 197412 211200
rect 443184 211080 443236 211132
rect 448520 211080 448572 211132
rect 516416 211080 516468 211132
rect 518348 211080 518400 211132
rect 442172 211012 442224 211064
rect 449164 211012 449216 211064
rect 370964 210264 371016 210316
rect 372712 210264 372764 210316
rect 373264 210264 373316 210316
rect 182916 209788 182968 209840
rect 197360 209788 197412 209840
rect 516140 209516 516192 209568
rect 519176 209516 519228 209568
rect 370964 209176 371016 209228
rect 372896 209176 372948 209228
rect 445668 209108 445720 209160
rect 450544 209108 450596 209160
rect 461584 209108 461636 209160
rect 303068 209040 303120 209092
rect 303528 209040 303580 209092
rect 342904 209040 342956 209092
rect 444564 209040 444616 209092
rect 445116 209040 445168 209092
rect 464344 209040 464396 209092
rect 372896 208360 372948 208412
rect 373356 208360 373408 208412
rect 445116 208292 445168 208344
rect 449256 208292 449308 208344
rect 370964 208088 371016 208140
rect 374000 208088 374052 208140
rect 445668 207612 445720 207664
rect 454684 207612 454736 207664
rect 181628 207000 181680 207052
rect 197360 207000 197412 207052
rect 516140 206864 516192 206916
rect 528652 206864 528704 206916
rect 515404 206796 515456 206848
rect 580172 206796 580224 206848
rect 302240 206116 302292 206168
rect 304264 206116 304316 206168
rect 444380 205844 444432 205896
rect 448152 205844 448204 205896
rect 516140 205844 516192 205896
rect 517796 205844 517848 205896
rect 444288 205708 444340 205760
rect 444656 205708 444708 205760
rect 180248 205640 180300 205692
rect 197360 205640 197412 205692
rect 443644 205572 443696 205624
rect 444196 205572 444248 205624
rect 447968 205572 448020 205624
rect 442908 205300 442960 205352
rect 446680 205300 446732 205352
rect 516140 204892 516192 204944
rect 516324 204892 516376 204944
rect 525892 204892 525944 204944
rect 444380 204756 444432 204808
rect 447784 204756 447836 204808
rect 516140 204212 516192 204264
rect 524604 204212 524656 204264
rect 442724 203940 442776 203992
rect 446404 203940 446456 203992
rect 442356 203328 442408 203380
rect 446588 203328 446640 203380
rect 173256 202852 173308 202904
rect 198280 202852 198332 202904
rect 3424 202784 3476 202836
rect 28264 202784 28316 202836
rect 447232 202784 447284 202836
rect 447876 202784 447928 202836
rect 516140 202784 516192 202836
rect 521752 202784 521804 202836
rect 442908 202716 442960 202768
rect 446496 202716 446548 202768
rect 371608 202308 371660 202360
rect 371884 202308 371936 202360
rect 173164 201492 173216 201544
rect 197360 201492 197412 201544
rect 445668 201492 445720 201544
rect 447232 201492 447284 201544
rect 514668 201220 514720 201272
rect 520648 201220 520700 201272
rect 445208 200064 445260 200116
rect 445392 200064 445444 200116
rect 514208 200064 514260 200116
rect 525800 200064 525852 200116
rect 514116 199996 514168 200048
rect 523040 199996 523092 200048
rect 303436 199384 303488 199436
rect 346308 199384 346360 199436
rect 173440 198704 173492 198756
rect 197544 198704 197596 198756
rect 514116 198636 514168 198688
rect 520280 198636 520332 198688
rect 445300 198024 445352 198076
rect 513564 198024 513616 198076
rect 476488 197956 476540 198008
rect 513380 197956 513432 198008
rect 444932 197752 444984 197804
rect 445300 197752 445352 197804
rect 370964 197616 371016 197668
rect 372620 197616 372672 197668
rect 374092 197616 374144 197668
rect 173348 197344 173400 197396
rect 197360 197344 197412 197396
rect 369124 197344 369176 197396
rect 369308 197344 369360 197396
rect 445300 197344 445352 197396
rect 476488 197344 476540 197396
rect 476764 197344 476816 197396
rect 445760 197276 445812 197328
rect 369860 197208 369912 197260
rect 371148 197208 371200 197260
rect 443368 197208 443420 197260
rect 445392 197208 445444 197260
rect 447140 197208 447192 197260
rect 513288 197276 513340 197328
rect 514944 197276 514996 197328
rect 516508 197208 516560 197260
rect 445208 197140 445260 197192
rect 445484 197140 445536 197192
rect 516324 197140 516376 197192
rect 466920 196800 466972 196852
rect 514208 196800 514260 196852
rect 447140 196664 447192 196716
rect 457444 196664 457496 196716
rect 514116 196664 514168 196716
rect 302792 196596 302844 196648
rect 369860 196596 369912 196648
rect 445576 196596 445628 196648
rect 460204 196596 460256 196648
rect 516140 196596 516192 196648
rect 445760 196052 445812 196104
rect 446496 196052 446548 196104
rect 445668 195984 445720 196036
rect 466920 195984 466972 196036
rect 346308 195304 346360 195356
rect 381544 195304 381596 195356
rect 303344 195236 303396 195288
rect 370320 195236 370372 195288
rect 445944 195236 445996 195288
rect 173532 194556 173584 194608
rect 197544 194556 197596 194608
rect 305644 194488 305696 194540
rect 510896 194488 510948 194540
rect 359464 194420 359516 194472
rect 366916 194420 366968 194472
rect 371976 194420 372028 194472
rect 375380 194420 375432 194472
rect 443276 194420 443328 194472
rect 506848 194420 506900 194472
rect 507768 194420 507820 194472
rect 514760 194420 514812 194472
rect 508872 194352 508924 194404
rect 514852 194352 514904 194404
rect 305736 193808 305788 193860
rect 438952 193808 439004 193860
rect 173624 193196 173676 193248
rect 197360 193196 197412 193248
rect 302608 193196 302660 193248
rect 371056 193196 371108 193248
rect 371976 193196 372028 193248
rect 522304 193128 522356 193180
rect 580172 193128 580224 193180
rect 302424 191768 302476 191820
rect 369216 191768 369268 191820
rect 370964 191768 371016 191820
rect 371700 191768 371752 191820
rect 371700 191088 371752 191140
rect 442264 191088 442316 191140
rect 193956 190884 194008 190936
rect 198280 190884 198332 190936
rect 172428 190068 172480 190120
rect 175924 190068 175976 190120
rect 352564 189728 352616 189780
rect 374460 189728 374512 189780
rect 375288 189728 375340 189780
rect 176108 189048 176160 189100
rect 197360 189048 197412 189100
rect 375288 189048 375340 189100
rect 446404 189048 446456 189100
rect 3424 188980 3476 189032
rect 155224 188980 155276 189032
rect 172428 188980 172480 189032
rect 181444 188980 181496 189032
rect 172428 187620 172480 187672
rect 188344 187620 188396 187672
rect 376944 187620 376996 187672
rect 443460 187620 443512 187672
rect 303068 186940 303120 186992
rect 303436 186940 303488 186992
rect 376944 186940 376996 186992
rect 174728 186328 174780 186380
rect 197360 186328 197412 186380
rect 172428 186192 172480 186244
rect 180064 186192 180116 186244
rect 196808 184968 196860 185020
rect 198464 184968 198516 185020
rect 172336 184832 172388 184884
rect 193864 184832 193916 184884
rect 302792 184832 302844 184884
rect 376852 184832 376904 184884
rect 378048 184832 378100 184884
rect 172428 184764 172480 184816
rect 186964 184764 187016 184816
rect 378048 184152 378100 184204
rect 399484 184152 399536 184204
rect 442172 184152 442224 184204
rect 172428 183472 172480 183524
rect 184204 183472 184256 183524
rect 178868 182180 178920 182232
rect 197360 182180 197412 182232
rect 172428 182112 172480 182164
rect 182824 182112 182876 182164
rect 302700 182112 302752 182164
rect 377680 182112 377732 182164
rect 378048 182112 378100 182164
rect 378048 181432 378100 181484
rect 395344 181432 395396 181484
rect 443092 181432 443144 181484
rect 195428 180888 195480 180940
rect 198280 180888 198332 180940
rect 172428 180752 172480 180804
rect 181536 180752 181588 180804
rect 373632 179392 373684 179444
rect 303344 179324 303396 179376
rect 304908 179324 304960 179376
rect 536104 179324 536156 179376
rect 580172 179324 580224 179376
rect 171140 179188 171192 179240
rect 180156 179188 180208 179240
rect 373540 178644 373592 178696
rect 442264 178644 442316 178696
rect 180340 178032 180392 178084
rect 197360 178032 197412 178084
rect 172244 177964 172296 178016
rect 196624 177964 196676 178016
rect 172428 177896 172480 177948
rect 178776 177896 178828 177948
rect 188344 176672 188396 176724
rect 197360 176672 197412 176724
rect 172244 176604 172296 176656
rect 195244 176604 195296 176656
rect 368388 176604 368440 176656
rect 372804 176604 372856 176656
rect 441988 176604 442040 176656
rect 302240 175244 302292 175296
rect 357256 175244 357308 175296
rect 358084 175244 358136 175296
rect 441988 175244 442040 175296
rect 442356 175244 442408 175296
rect 172428 175176 172480 175228
rect 192576 175176 192628 175228
rect 186964 173884 187016 173936
rect 197728 173884 197780 173936
rect 172428 173816 172480 173868
rect 191196 173816 191248 173868
rect 184204 172524 184256 172576
rect 197360 172524 197412 172576
rect 372436 172524 372488 172576
rect 442724 172524 442776 172576
rect 444748 172524 444800 172576
rect 172428 172388 172480 172440
rect 177396 172388 177448 172440
rect 373448 171776 373500 171828
rect 442448 171776 442500 171828
rect 172428 171028 172480 171080
rect 198096 171028 198148 171080
rect 442632 171028 442684 171080
rect 445116 171028 445168 171080
rect 371240 170484 371292 170536
rect 371884 170484 371936 170536
rect 371240 170348 371292 170400
rect 376024 170348 376076 170400
rect 442632 170348 442684 170400
rect 172244 169668 172296 169720
rect 195336 169668 195388 169720
rect 371700 169260 371752 169312
rect 372436 169260 372488 169312
rect 302792 168988 302844 169040
rect 371700 168988 371752 169040
rect 373724 168308 373776 168360
rect 374368 168308 374420 168360
rect 441804 168308 441856 168360
rect 445116 168308 445168 168360
rect 178776 167628 178828 167680
rect 197452 167628 197504 167680
rect 371884 167628 371936 167680
rect 444840 167628 444892 167680
rect 444840 167288 444892 167340
rect 445024 167288 445076 167340
rect 182824 167016 182876 167068
rect 197360 167016 197412 167068
rect 172428 166948 172480 167000
rect 196716 166948 196768 167000
rect 301504 166948 301556 167000
rect 580172 166948 580224 167000
rect 302792 166268 302844 166320
rect 371976 166268 372028 166320
rect 372344 166268 372396 166320
rect 172152 165520 172204 165572
rect 174636 165520 174688 165572
rect 373356 165520 373408 165572
rect 441896 165520 441948 165572
rect 443000 165520 443052 165572
rect 3240 164160 3292 164212
rect 11704 164160 11756 164212
rect 172244 164160 172296 164212
rect 198740 164160 198792 164212
rect 369032 164160 369084 164212
rect 371240 164160 371292 164212
rect 444656 163752 444708 163804
rect 445300 163752 445352 163804
rect 171784 163616 171836 163668
rect 180340 163616 180392 163668
rect 371976 163480 372028 163532
rect 372344 163480 372396 163532
rect 444656 163480 444708 163532
rect 180064 162868 180116 162920
rect 197544 162868 197596 162920
rect 302792 162868 302844 162920
rect 369032 162868 369084 162920
rect 442908 162800 442960 162852
rect 445208 162800 445260 162852
rect 181444 162120 181496 162172
rect 198464 162120 198516 162172
rect 372252 161440 372304 161492
rect 442908 161440 442960 161492
rect 172428 161236 172480 161288
rect 176016 161236 176068 161288
rect 445852 160828 445904 160880
rect 446496 160828 446548 160880
rect 169208 160692 169260 160744
rect 178684 160692 178736 160744
rect 373264 160692 373316 160744
rect 445852 160692 445904 160744
rect 177396 158720 177448 158772
rect 197544 158720 197596 158772
rect 302516 158720 302568 158772
rect 166908 158652 166960 158704
rect 170404 158652 170456 158704
rect 374184 158652 374236 158704
rect 164884 158584 164936 158636
rect 170496 158584 170548 158636
rect 162860 158516 162912 158568
rect 174544 158516 174596 158568
rect 302884 157972 302936 158024
rect 369400 157972 369452 158024
rect 374184 157972 374236 158024
rect 443092 157972 443144 158024
rect 443644 157972 443696 158024
rect 175924 157360 175976 157412
rect 197360 157360 197412 157412
rect 171968 156612 172020 156664
rect 188344 156612 188396 156664
rect 369860 156612 369912 156664
rect 374276 156612 374328 156664
rect 445208 156612 445260 156664
rect 393964 156476 394016 156528
rect 394608 156476 394660 156528
rect 394608 156204 394660 156256
rect 513380 156204 513432 156256
rect 370504 156136 370556 156188
rect 371056 156136 371108 156188
rect 515036 156136 515088 156188
rect 370596 156068 370648 156120
rect 371148 156068 371200 156120
rect 515128 156068 515180 156120
rect 370136 156000 370188 156052
rect 370964 156000 371016 156052
rect 515312 156000 515364 156052
rect 369400 155932 369452 155984
rect 516968 155932 517020 155984
rect 302976 155184 303028 155236
rect 370228 155184 370280 155236
rect 374644 155184 374696 155236
rect 441620 155320 441672 155372
rect 507768 155252 507820 155304
rect 514024 155252 514076 155304
rect 468484 155184 468536 155236
rect 516600 155184 516652 155236
rect 370228 154640 370280 154692
rect 174544 154572 174596 154624
rect 197544 154572 197596 154624
rect 515220 154572 515272 154624
rect 172336 154504 172388 154556
rect 188436 154504 188488 154556
rect 368388 154504 368440 154556
rect 369676 154504 369728 154556
rect 373632 154504 373684 154556
rect 441804 154504 441856 154556
rect 444564 154504 444616 154556
rect 444748 154504 444800 154556
rect 445208 154504 445260 154556
rect 459744 154504 459796 154556
rect 460204 154504 460256 154556
rect 172244 154436 172296 154488
rect 187056 154436 187108 154488
rect 442448 154436 442500 154488
rect 445576 154436 445628 154488
rect 442356 154368 442408 154420
rect 444656 154368 444708 154420
rect 441620 154300 441672 154352
rect 444840 154300 444892 154352
rect 437388 154164 437440 154216
rect 441712 154164 441764 154216
rect 489184 154164 489236 154216
rect 514116 154164 514168 154216
rect 485044 154096 485096 154148
rect 513656 154096 513708 154148
rect 482284 154028 482336 154080
rect 513748 154028 513800 154080
rect 359648 153960 359700 154012
rect 368388 153960 368440 154012
rect 459744 153960 459796 154012
rect 513196 153960 513248 154012
rect 302792 153892 302844 153944
rect 370044 153892 370096 153944
rect 446404 153892 446456 153944
rect 516784 153892 516836 153944
rect 303528 153824 303580 153876
rect 372620 153824 372672 153876
rect 431868 153824 431920 153876
rect 434720 153824 434772 153876
rect 444748 153824 444800 153876
rect 515404 153824 515456 153876
rect 445300 153756 445352 153808
rect 514392 153756 514444 153808
rect 445116 153688 445168 153740
rect 514576 153688 514628 153740
rect 444656 153620 444708 153672
rect 513840 153620 513892 153672
rect 444840 153552 444892 153604
rect 514484 153552 514536 153604
rect 442264 153484 442316 153536
rect 514208 153484 514260 153536
rect 445576 153416 445628 153468
rect 514300 153416 514352 153468
rect 443092 153348 443144 153400
rect 514760 153348 514812 153400
rect 359004 153280 359056 153332
rect 188344 153212 188396 153264
rect 197360 153212 197412 153264
rect 302700 153212 302752 153264
rect 369860 153212 369912 153264
rect 172428 153144 172480 153196
rect 184296 153144 184348 153196
rect 369216 153144 369268 153196
rect 372436 153144 372488 153196
rect 431316 153280 431368 153332
rect 514668 153280 514720 153332
rect 372620 153212 372672 153264
rect 372988 153212 373040 153264
rect 515588 153212 515640 153264
rect 373724 153144 373776 153196
rect 479524 153144 479576 153196
rect 513288 153144 513340 153196
rect 520924 153144 520976 153196
rect 580172 153144 580224 153196
rect 172336 153076 172388 153128
rect 182916 153076 182968 153128
rect 370044 153076 370096 153128
rect 372620 153076 372672 153128
rect 373540 153076 373592 153128
rect 493324 153076 493376 153128
rect 513472 153076 513524 153128
rect 516232 153076 516284 153128
rect 528836 153076 528888 153128
rect 342168 153008 342220 153060
rect 371240 153008 371292 153060
rect 516140 153008 516192 153060
rect 518900 153008 518952 153060
rect 357348 152940 357400 152992
rect 369492 152940 369544 152992
rect 307668 152872 307720 152924
rect 369584 152872 369636 152924
rect 497464 152872 497516 152924
rect 516692 152872 516744 152924
rect 313188 152804 313240 152856
rect 369308 152804 369360 152856
rect 494704 152804 494756 152856
rect 516508 152804 516560 152856
rect 357256 152736 357308 152788
rect 372712 152736 372764 152788
rect 490564 152736 490616 152788
rect 513380 152736 513432 152788
rect 340788 152668 340840 152720
rect 371240 152668 371292 152720
rect 475384 152668 475436 152720
rect 516324 152668 516376 152720
rect 303068 152600 303120 152652
rect 369216 152600 369268 152652
rect 472624 152600 472676 152652
rect 302792 152532 302844 152584
rect 370044 152532 370096 152584
rect 374644 152532 374696 152584
rect 471244 152532 471296 152584
rect 303436 152464 303488 152516
rect 372896 152464 372948 152516
rect 445668 152464 445720 152516
rect 450544 152464 450596 152516
rect 516140 152532 516192 152584
rect 516416 152464 516468 152516
rect 513932 152124 513984 152176
rect 442724 152056 442776 152108
rect 514944 152056 514996 152108
rect 372712 151988 372764 152040
rect 441804 151988 441856 152040
rect 444748 151988 444800 152040
rect 514852 151988 514904 152040
rect 431408 151920 431460 151972
rect 513104 151920 513156 151972
rect 516508 151920 516560 151972
rect 359556 151852 359608 151904
rect 372896 151852 372948 151904
rect 515496 151852 515548 151904
rect 516324 151852 516376 151904
rect 442632 151784 442684 151836
rect 444196 151784 444248 151836
rect 516508 151784 516560 151836
rect 516968 151784 517020 151836
rect 171692 151716 171744 151768
rect 181628 151716 181680 151768
rect 302792 151716 302844 151768
rect 359004 151716 359056 151768
rect 369768 151716 369820 151768
rect 373448 151716 373500 151768
rect 514116 151716 514168 151768
rect 444380 151648 444432 151700
rect 444748 151648 444800 151700
rect 514208 151648 514260 151700
rect 513564 151580 513616 151632
rect 514392 151648 514444 151700
rect 171508 151444 171560 151496
rect 180248 151444 180300 151496
rect 514300 151444 514352 151496
rect 514300 150628 514352 150680
rect 171600 150560 171652 150612
rect 173256 150560 173308 150612
rect 187056 150424 187108 150476
rect 197544 150424 197596 150476
rect 3424 150356 3476 150408
rect 29644 150356 29696 150408
rect 171692 150356 171744 150408
rect 173164 150356 173216 150408
rect 171692 149404 171744 149456
rect 173440 149404 173492 149456
rect 184296 149064 184348 149116
rect 197360 149064 197412 149116
rect 172244 148860 172296 148912
rect 173348 148860 173400 148912
rect 171692 148792 171744 148844
rect 173532 148792 173584 148844
rect 173164 148316 173216 148368
rect 198096 148316 198148 148368
rect 371332 148248 371384 148300
rect 375472 148248 375524 148300
rect 171508 147840 171560 147892
rect 173624 147840 173676 147892
rect 172428 147568 172480 147620
rect 193956 147568 194008 147620
rect 171508 147500 171560 147552
rect 176108 147500 176160 147552
rect 371332 147228 371384 147280
rect 375564 147228 375616 147280
rect 513380 147092 513432 147144
rect 513564 147092 513616 147144
rect 513656 147024 513708 147076
rect 514484 147024 514536 147076
rect 513564 146956 513616 147008
rect 514392 146956 514444 147008
rect 513748 146888 513800 146940
rect 514576 146888 514628 146940
rect 369216 146820 369268 146872
rect 369768 146820 369820 146872
rect 371976 146820 372028 146872
rect 375656 146820 375708 146872
rect 372620 146752 372672 146804
rect 373724 146752 373776 146804
rect 182916 146276 182968 146328
rect 197636 146276 197688 146328
rect 172428 146208 172480 146260
rect 196808 146208 196860 146260
rect 371976 146208 372028 146260
rect 393964 146208 394016 146260
rect 172336 146140 172388 146192
rect 174728 146140 174780 146192
rect 171508 145800 171560 145852
rect 178868 145800 178920 145852
rect 371332 145596 371384 145648
rect 375932 145596 375984 145648
rect 371332 145460 371384 145512
rect 375840 145460 375892 145512
rect 181536 144916 181588 144968
rect 197360 144916 197412 144968
rect 172428 144848 172480 144900
rect 195428 144848 195480 144900
rect 302792 144848 302844 144900
rect 359648 144848 359700 144900
rect 515404 144848 515456 144900
rect 516140 144848 516192 144900
rect 371332 144508 371384 144560
rect 375748 144508 375800 144560
rect 171600 144168 171652 144220
rect 184204 144168 184256 144220
rect 371332 144100 371384 144152
rect 374460 144100 374512 144152
rect 172244 143488 172296 143540
rect 186964 143488 187016 143540
rect 371332 143420 371384 143472
rect 406384 143488 406436 143540
rect 431408 143488 431460 143540
rect 371976 143012 372028 143064
rect 372988 143012 373040 143064
rect 171508 142808 171560 142860
rect 182824 142808 182876 142860
rect 179420 142128 179472 142180
rect 197360 142128 197412 142180
rect 172428 142060 172480 142112
rect 181444 142060 181496 142112
rect 302332 142060 302384 142112
rect 359556 142060 359608 142112
rect 371976 142060 372028 142112
rect 381544 142060 381596 142112
rect 431316 142060 431368 142112
rect 171416 141924 171468 141976
rect 178776 141924 178828 141976
rect 171508 141244 171560 141296
rect 180064 141244 180116 141296
rect 178040 140768 178092 140820
rect 197360 140768 197412 140820
rect 372620 140360 372672 140412
rect 372988 140360 373040 140412
rect 172244 140020 172296 140072
rect 187056 140020 187108 140072
rect 171692 139748 171744 139800
rect 173164 139748 173216 139800
rect 371700 139340 371752 139392
rect 371976 139340 372028 139392
rect 372160 139340 372212 139392
rect 372896 139340 372948 139392
rect 518164 139340 518216 139392
rect 580172 139340 580224 139392
rect 172428 139272 172480 139324
rect 177396 139272 177448 139324
rect 371332 139272 371384 139324
rect 395344 139272 395396 139324
rect 395988 139272 396040 139324
rect 371700 139204 371752 139256
rect 399484 139204 399536 139256
rect 171876 138864 171928 138916
rect 175924 138864 175976 138916
rect 171692 138728 171744 138780
rect 174544 138728 174596 138780
rect 399484 138728 399536 138780
rect 431316 138728 431368 138780
rect 395988 138660 396040 138712
rect 429844 138660 429896 138712
rect 175924 137980 175976 138032
rect 197360 137980 197412 138032
rect 445852 137980 445904 138032
rect 446404 137980 446456 138032
rect 3240 137912 3292 137964
rect 152464 137912 152516 137964
rect 172428 137912 172480 137964
rect 188344 137912 188396 137964
rect 371332 137572 371384 137624
rect 373632 137572 373684 137624
rect 371332 137300 371384 137352
rect 371516 137300 371568 137352
rect 172336 137232 172388 137284
rect 184296 137232 184348 137284
rect 172520 136620 172572 136672
rect 197360 136620 197412 136672
rect 445300 136620 445352 136672
rect 497464 136620 497516 136672
rect 172428 136552 172480 136604
rect 182916 136552 182968 136604
rect 172244 136484 172296 136536
rect 181536 136484 181588 136536
rect 170404 135872 170456 135924
rect 198004 135872 198056 135924
rect 441620 135872 441672 135924
rect 447232 135872 447284 135924
rect 500224 135872 500276 135924
rect 172244 135260 172296 135312
rect 179420 135260 179472 135312
rect 445024 135260 445076 135312
rect 445668 135260 445720 135312
rect 503076 135260 503128 135312
rect 171692 135192 171744 135244
rect 175924 135192 175976 135244
rect 369124 135192 369176 135244
rect 171876 135124 171928 135176
rect 178040 135124 178092 135176
rect 369124 134852 369176 134904
rect 371700 134308 371752 134360
rect 374184 134308 374236 134360
rect 443092 133968 443144 134020
rect 490564 133968 490616 134020
rect 172428 133900 172480 133952
rect 197728 133900 197780 133952
rect 442908 133900 442960 133952
rect 445116 133900 445168 133952
rect 503168 133900 503220 133952
rect 371516 132948 371568 133000
rect 372988 132948 373040 133000
rect 171140 132472 171192 132524
rect 197360 132472 197412 132524
rect 442816 132472 442868 132524
rect 444196 132472 444248 132524
rect 445116 132472 445168 132524
rect 503260 132472 503312 132524
rect 172428 131044 172480 131096
rect 197360 131044 197412 131096
rect 370044 130432 370096 130484
rect 373264 130432 373316 130484
rect 370320 130364 370372 130416
rect 373356 130364 373408 130416
rect 172244 129956 172296 130008
rect 178040 129956 178092 130008
rect 444840 129004 444892 129056
rect 476764 129004 476816 129056
rect 503628 129004 503680 129056
rect 172336 128256 172388 128308
rect 197360 128256 197412 128308
rect 442908 127644 442960 127696
rect 504272 127644 504324 127696
rect 443368 127576 443420 127628
rect 444932 127576 444984 127628
rect 504364 127576 504416 127628
rect 171324 126896 171376 126948
rect 197636 126896 197688 126948
rect 526444 126896 526496 126948
rect 580172 126896 580224 126948
rect 444932 126284 444984 126336
rect 467104 126284 467156 126336
rect 493968 126284 494020 126336
rect 444840 126216 444892 126268
rect 457444 126216 457496 126268
rect 494704 126216 494756 126268
rect 371608 126012 371660 126064
rect 441896 126012 441948 126064
rect 371700 125944 371752 125996
rect 442908 125944 442960 125996
rect 370412 125876 370464 125928
rect 371332 125876 371384 125928
rect 443368 125876 443420 125928
rect 172244 125740 172296 125792
rect 180064 125740 180116 125792
rect 172428 125672 172480 125724
rect 181444 125672 181496 125724
rect 172336 125604 172388 125656
rect 182824 125604 182876 125656
rect 371424 125468 371476 125520
rect 441804 125468 441856 125520
rect 444932 125468 444984 125520
rect 369308 125400 369360 125452
rect 443092 125400 443144 125452
rect 374828 125332 374880 125384
rect 442080 125332 442132 125384
rect 444840 125332 444892 125384
rect 302424 125196 302476 125248
rect 369952 125196 370004 125248
rect 302516 125128 302568 125180
rect 369860 125128 369912 125180
rect 441620 125264 441672 125316
rect 302884 125060 302936 125112
rect 370044 125060 370096 125112
rect 302700 124992 302752 125044
rect 369308 124992 369360 125044
rect 302976 124924 303028 124976
rect 370320 124924 370372 124976
rect 445760 125196 445812 125248
rect 513196 125196 513248 125248
rect 493968 125128 494020 125180
rect 513380 125128 513432 125180
rect 494704 125060 494756 125112
rect 500224 124992 500276 125044
rect 513288 124992 513340 125044
rect 513380 124992 513432 125044
rect 446404 124924 446456 124976
rect 516140 124924 516192 124976
rect 172520 124856 172572 124908
rect 197452 124856 197504 124908
rect 302240 124856 302292 124908
rect 370228 124856 370280 124908
rect 370872 124856 370924 124908
rect 441620 124856 441672 124908
rect 490564 124856 490616 124908
rect 513472 124856 513524 124908
rect 497464 124788 497516 124840
rect 516232 124788 516284 124840
rect 369860 124720 369912 124772
rect 374092 124720 374144 124772
rect 374828 124720 374880 124772
rect 429844 124720 429896 124772
rect 516324 124720 516376 124772
rect 171508 124312 171560 124364
rect 175924 124312 175976 124364
rect 171876 124244 171928 124296
rect 174544 124244 174596 124296
rect 172152 124176 172204 124228
rect 173164 124176 173216 124228
rect 178040 124108 178092 124160
rect 197360 124108 197412 124160
rect 431316 124108 431368 124160
rect 516508 124108 516560 124160
rect 368204 124040 368256 124092
rect 369400 124040 369452 124092
rect 503076 124040 503128 124092
rect 513840 124040 513892 124092
rect 503168 123972 503220 124024
rect 513748 123972 513800 124024
rect 503628 123904 503680 123956
rect 513564 123904 513616 123956
rect 503260 123836 503312 123888
rect 513932 123836 513984 123888
rect 504364 123768 504416 123820
rect 513656 123768 513708 123820
rect 504272 123700 504324 123752
rect 514116 123700 514168 123752
rect 302976 123496 303028 123548
rect 370412 123496 370464 123548
rect 302884 123428 302936 123480
rect 369860 123428 369912 123480
rect 168932 122884 168984 122936
rect 177304 122884 177356 122936
rect 160928 122816 160980 122868
rect 192484 122816 192536 122868
rect 320824 122816 320876 122868
rect 510896 122816 510948 122868
rect 164884 122748 164936 122800
rect 170404 122748 170456 122800
rect 162860 122680 162912 122732
rect 191104 122748 191156 122800
rect 431868 122748 431920 122800
rect 434720 122748 434772 122800
rect 441252 122748 441304 122800
rect 512920 122748 512972 122800
rect 433156 122680 433208 122732
rect 504916 122680 504968 122732
rect 506848 122680 506900 122732
rect 514024 122680 514076 122732
rect 437204 122612 437256 122664
rect 441712 122612 441764 122664
rect 508872 122612 508924 122664
rect 309784 122544 309836 122596
rect 438860 122544 438912 122596
rect 301504 122068 301556 122120
rect 366916 122068 366968 122120
rect 172060 120028 172112 120080
rect 197360 120028 197412 120080
rect 302516 120028 302568 120080
rect 370136 120028 370188 120080
rect 171876 118600 171928 118652
rect 197636 118600 197688 118652
rect 302608 117240 302660 117292
rect 368204 117240 368256 117292
rect 171968 115880 172020 115932
rect 198556 115880 198608 115932
rect 171784 114452 171836 114504
rect 197544 114452 197596 114504
rect 318064 113092 318116 113144
rect 579804 113092 579856 113144
rect 175924 112412 175976 112464
rect 197452 112412 197504 112464
rect 3424 111732 3476 111784
rect 159364 111732 159416 111784
rect 182824 111732 182876 111784
rect 197360 111732 197412 111784
rect 302516 111732 302568 111784
rect 370504 111732 370556 111784
rect 181444 110372 181496 110424
rect 197544 110372 197596 110424
rect 302792 108944 302844 108996
rect 371424 108944 371476 108996
rect 180064 107584 180116 107636
rect 198004 107584 198056 107636
rect 174544 103436 174596 103488
rect 198004 103436 198056 103488
rect 173164 102076 173216 102128
rect 198004 102076 198056 102128
rect 302792 102076 302844 102128
rect 369860 102076 369912 102128
rect 533344 100648 533396 100700
rect 580172 100648 580224 100700
rect 232044 99968 232096 100020
rect 232320 99900 232372 99952
rect 298928 99696 298980 99748
rect 322204 99696 322256 99748
rect 299112 99628 299164 99680
rect 323584 99628 323636 99680
rect 298652 99560 298704 99612
rect 359464 99560 359516 99612
rect 299480 99492 299532 99544
rect 431224 99492 431276 99544
rect 211620 99424 211672 99476
rect 211804 99424 211856 99476
rect 299848 99424 299900 99476
rect 501604 99424 501656 99476
rect 166908 99356 166960 99408
rect 298284 99356 298336 99408
rect 299664 99356 299716 99408
rect 502984 99356 503036 99408
rect 298468 99288 298520 99340
rect 301504 99288 301556 99340
rect 101404 99220 101456 99272
rect 211988 99220 212040 99272
rect 299296 99220 299348 99272
rect 305736 99288 305788 99340
rect 94504 99152 94556 99204
rect 207848 99152 207900 99204
rect 271420 99152 271472 99204
rect 423772 99152 423824 99204
rect 93124 99084 93176 99136
rect 213828 99084 213880 99136
rect 273812 99084 273864 99136
rect 435364 99084 435416 99136
rect 71044 99016 71096 99068
rect 210240 99016 210292 99068
rect 275008 99016 275060 99068
rect 440884 99016 440936 99068
rect 57244 98948 57296 99000
rect 207664 98948 207716 99000
rect 290096 98948 290148 99000
rect 457444 98948 457496 99000
rect 50344 98880 50396 98932
rect 207020 98880 207072 98932
rect 277400 98880 277452 98932
rect 458180 98880 458232 98932
rect 46204 98812 46256 98864
rect 205824 98812 205876 98864
rect 279148 98812 279200 98864
rect 467104 98812 467156 98864
rect 36544 98744 36596 98796
rect 202236 98744 202288 98796
rect 282920 98744 282972 98796
rect 490564 98744 490616 98796
rect 29644 98676 29696 98728
rect 204628 98676 204680 98728
rect 292948 98676 293000 98728
rect 550640 98676 550692 98728
rect 19248 98608 19300 98660
rect 203064 98608 203116 98660
rect 293500 98608 293552 98660
rect 554780 98608 554832 98660
rect 263048 98540 263100 98592
rect 374000 98540 374052 98592
rect 258632 98472 258684 98524
rect 345664 98472 345716 98524
rect 256884 98404 256936 98456
rect 336004 98404 336056 98456
rect 218520 98336 218572 98388
rect 218980 98336 219032 98388
rect 270776 98336 270828 98388
rect 413284 98336 413336 98388
rect 201592 98268 201644 98320
rect 201868 98268 201920 98320
rect 208492 98268 208544 98320
rect 208860 98268 208912 98320
rect 270960 98268 271012 98320
rect 414664 98268 414716 98320
rect 289360 98200 289412 98252
rect 289636 98200 289688 98252
rect 150348 97928 150400 97980
rect 225144 97928 225196 97980
rect 238116 97928 238168 97980
rect 238760 97928 238812 97980
rect 134524 97860 134576 97912
rect 214380 97860 214432 97912
rect 215300 97860 215352 97912
rect 222384 97860 222436 97912
rect 238024 97860 238076 97912
rect 239680 97860 239732 97912
rect 126888 97792 126940 97844
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 124864 97724 124916 97776
rect 215116 97792 215168 97844
rect 219808 97792 219860 97844
rect 234620 97792 234672 97844
rect 239312 97792 239364 97844
rect 251640 97792 251692 97844
rect 256700 97792 256752 97844
rect 264612 97792 264664 97844
rect 322204 97928 322256 97980
rect 272708 97860 272760 97912
rect 327724 97860 327776 97912
rect 126244 97656 126296 97708
rect 208952 97656 209004 97708
rect 216680 97724 216732 97776
rect 226340 97724 226392 97776
rect 242072 97724 242124 97776
rect 253296 97724 253348 97776
rect 259276 97724 259328 97776
rect 267280 97724 267332 97776
rect 268200 97724 268252 97776
rect 276020 97792 276072 97844
rect 278136 97792 278188 97844
rect 352564 97792 352616 97844
rect 275376 97724 275428 97776
rect 282184 97724 282236 97776
rect 282736 97724 282788 97776
rect 359464 97724 359516 97776
rect 119344 97588 119396 97640
rect 221188 97656 221240 97708
rect 227720 97656 227772 97708
rect 229560 97656 229612 97708
rect 247316 97656 247368 97708
rect 253204 97656 253256 97708
rect 254032 97656 254084 97708
rect 262772 97656 262824 97708
rect 262956 97656 263008 97708
rect 267648 97656 267700 97708
rect 270592 97656 270644 97708
rect 115204 97520 115256 97572
rect 205732 97520 205784 97572
rect 216772 97588 216824 97640
rect 250444 97588 250496 97640
rect 262864 97588 262916 97640
rect 265808 97588 265860 97640
rect 272708 97588 272760 97640
rect 272984 97656 273036 97708
rect 277308 97588 277360 97640
rect 277768 97588 277820 97640
rect 282000 97588 282052 97640
rect 282276 97656 282328 97708
rect 363604 97656 363656 97708
rect 370504 97588 370556 97640
rect 218612 97520 218664 97572
rect 218796 97520 218848 97572
rect 224960 97520 225012 97572
rect 247500 97520 247552 97572
rect 258724 97520 258776 97572
rect 262588 97520 262640 97572
rect 369124 97520 369176 97572
rect 200212 97452 200264 97504
rect 200948 97452 201000 97504
rect 203340 97452 203392 97504
rect 206652 97452 206704 97504
rect 212540 97452 212592 97504
rect 224224 97452 224276 97504
rect 257436 97452 257488 97504
rect 263048 97452 263100 97504
rect 267740 97452 267792 97504
rect 273260 97452 273312 97504
rect 278964 97452 279016 97504
rect 282000 97452 282052 97504
rect 282184 97452 282236 97504
rect 425704 97452 425756 97504
rect 97264 97384 97316 97436
rect 58624 97316 58676 97368
rect 206008 97316 206060 97368
rect 215576 97384 215628 97436
rect 218060 97384 218112 97436
rect 232504 97384 232556 97436
rect 244464 97384 244516 97436
rect 248420 97384 248472 97436
rect 208124 97316 208176 97368
rect 227812 97316 227864 97368
rect 243268 97316 243320 97368
rect 256976 97384 257028 97436
rect 263416 97384 263468 97436
rect 271328 97384 271380 97436
rect 276572 97384 276624 97436
rect 429844 97384 429896 97436
rect 253296 97316 253348 97368
rect 258356 97316 258408 97368
rect 260472 97316 260524 97368
rect 276664 97316 276716 97368
rect 276756 97316 276808 97368
rect 277124 97316 277176 97368
rect 39948 97248 40000 97300
rect 203340 97248 203392 97300
rect 206928 97248 206980 97300
rect 227168 97248 227220 97300
rect 227628 97248 227680 97300
rect 238300 97248 238352 97300
rect 246304 97248 246356 97300
rect 271052 97248 271104 97300
rect 272432 97248 272484 97300
rect 282276 97316 282328 97368
rect 281080 97248 281132 97300
rect 281356 97248 281408 97300
rect 282000 97248 282052 97300
rect 285128 97248 285180 97300
rect 285588 97248 285640 97300
rect 285864 97316 285916 97368
rect 436744 97316 436796 97368
rect 443644 97248 443696 97300
rect 142804 97180 142856 97232
rect 208860 97180 208912 97232
rect 208952 97180 209004 97232
rect 221004 97180 221056 97232
rect 248420 97180 248472 97232
rect 260104 97180 260156 97232
rect 267280 97180 267332 97232
rect 196624 97112 196676 97164
rect 217968 97112 218020 97164
rect 219716 97112 219768 97164
rect 220360 97112 220412 97164
rect 231860 97112 231912 97164
rect 237748 97112 237800 97164
rect 240048 97112 240100 97164
rect 242716 97112 242768 97164
rect 261024 97112 261076 97164
rect 268844 97180 268896 97232
rect 269028 97180 269080 97232
rect 270040 97180 270092 97232
rect 271144 97180 271196 97232
rect 274180 97180 274232 97232
rect 274548 97180 274600 97232
rect 275560 97180 275612 97232
rect 275928 97180 275980 97232
rect 276020 97180 276072 97232
rect 323584 97180 323636 97232
rect 192484 97044 192536 97096
rect 202696 97044 202748 97096
rect 202788 97044 202840 97096
rect 205456 97044 205508 97096
rect 205732 97044 205784 97096
rect 219164 97044 219216 97096
rect 241336 97044 241388 97096
rect 242164 97044 242216 97096
rect 246672 97044 246724 97096
rect 246856 97044 246908 97096
rect 253480 97044 253532 97096
rect 253756 97044 253808 97096
rect 255044 97044 255096 97096
rect 198004 96976 198056 97028
rect 195244 96908 195296 96960
rect 201868 96908 201920 96960
rect 201960 96908 202012 96960
rect 202512 96908 202564 96960
rect 211436 96976 211488 97028
rect 241704 96976 241756 97028
rect 242532 96976 242584 97028
rect 250076 96976 250128 97028
rect 250720 96976 250772 97028
rect 251272 96976 251324 97028
rect 252192 96976 252244 97028
rect 252284 96976 252336 97028
rect 252468 96976 252520 97028
rect 254676 96976 254728 97028
rect 255136 96976 255188 97028
rect 208860 96908 208912 96960
rect 212632 96908 212684 96960
rect 215760 96908 215812 96960
rect 216312 96908 216364 96960
rect 216864 96908 216916 96960
rect 217140 96908 217192 96960
rect 219716 96908 219768 96960
rect 220452 96908 220504 96960
rect 221464 96908 221516 96960
rect 221924 96908 221976 96960
rect 222292 96908 222344 96960
rect 222936 96908 222988 96960
rect 234712 96908 234764 96960
rect 235448 96908 235500 96960
rect 236460 96908 236512 96960
rect 237196 96908 237248 96960
rect 237656 96908 237708 96960
rect 238392 96908 238444 96960
rect 239036 96908 239088 96960
rect 239404 96908 239456 96960
rect 240324 96908 240376 96960
rect 240784 96908 240836 96960
rect 241520 96908 241572 96960
rect 242440 96908 242492 96960
rect 243728 96908 243780 96960
rect 244096 96908 244148 96960
rect 244740 96908 244792 96960
rect 245384 96908 245436 96960
rect 245936 96908 245988 96960
rect 246580 96908 246632 96960
rect 247132 96908 247184 96960
rect 248236 96908 248288 96960
rect 248512 96908 248564 96960
rect 249340 96908 249392 96960
rect 250628 96908 250680 96960
rect 250996 96908 251048 96960
rect 251456 96908 251508 96960
rect 252008 96908 252060 96960
rect 252652 96908 252704 96960
rect 253664 96908 253716 96960
rect 254216 96908 254268 96960
rect 255044 96908 255096 96960
rect 199384 96840 199436 96892
rect 202788 96840 202840 96892
rect 203524 96840 203576 96892
rect 207204 96840 207256 96892
rect 222476 96840 222528 96892
rect 223304 96840 223356 96892
rect 234620 96840 234672 96892
rect 235816 96840 235868 96892
rect 240232 96840 240284 96892
rect 240968 96840 241020 96892
rect 242348 96840 242400 96892
rect 242808 96840 242860 96892
rect 245108 96840 245160 96892
rect 245476 96840 245528 96892
rect 246120 96840 246172 96892
rect 246948 96840 247000 96892
rect 248696 96840 248748 96892
rect 249524 96840 249576 96892
rect 250260 96840 250312 96892
rect 250812 96840 250864 96892
rect 251824 96840 251876 96892
rect 252284 96840 252336 96892
rect 265900 97044 265952 97096
rect 266176 97044 266228 97096
rect 298008 97112 298060 97164
rect 256056 96976 256108 97028
rect 256424 96976 256476 97028
rect 257252 96976 257304 97028
rect 257896 96976 257948 97028
rect 258080 96976 258132 97028
rect 259092 96976 259144 97028
rect 261760 96976 261812 97028
rect 262036 96976 262088 97028
rect 263600 96976 263652 97028
rect 264796 96976 264848 97028
rect 265440 96976 265492 97028
rect 267004 96976 267056 97028
rect 267188 97044 267240 97096
rect 267556 97044 267608 97096
rect 267648 97044 267700 97096
rect 302884 97112 302936 97164
rect 300124 96976 300176 97028
rect 255688 96908 255740 96960
rect 256148 96908 256200 96960
rect 256332 96908 256384 96960
rect 256608 96908 256660 96960
rect 257620 96908 257672 96960
rect 257988 96908 258040 96960
rect 258448 96908 258500 96960
rect 259000 96908 259052 96960
rect 259460 96908 259512 96960
rect 260288 96908 260340 96960
rect 261208 96908 261260 96960
rect 261852 96908 261904 96960
rect 264060 96908 264112 96960
rect 264520 96908 264572 96960
rect 265256 96908 265308 96960
rect 265992 96908 266044 96960
rect 266820 96908 266872 96960
rect 267372 96908 267424 96960
rect 268016 96908 268068 96960
rect 268660 96908 268712 96960
rect 269764 96908 269816 96960
rect 270224 96908 270276 96960
rect 271236 96908 271288 96960
rect 271788 96908 271840 96960
rect 272616 96908 272668 96960
rect 272892 96908 272944 96960
rect 273260 96908 273312 96960
rect 298836 96908 298888 96960
rect 98644 96772 98696 96824
rect 204076 96772 204128 96824
rect 215484 96772 215536 96824
rect 216496 96772 216548 96824
rect 217140 96772 217192 96824
rect 217692 96772 217744 96824
rect 218244 96772 218296 96824
rect 218888 96772 218940 96824
rect 219440 96772 219492 96824
rect 220452 96772 220504 96824
rect 221096 96772 221148 96824
rect 221648 96772 221700 96824
rect 222292 96772 222344 96824
rect 223120 96772 223172 96824
rect 231584 96772 231636 96824
rect 237104 96772 237156 96824
rect 240692 96772 240744 96824
rect 241336 96772 241388 96824
rect 241888 96772 241940 96824
rect 242716 96772 242768 96824
rect 245660 96772 245712 96824
rect 246764 96772 246816 96824
rect 253388 96772 253440 96824
rect 253848 96772 253900 96824
rect 254768 96772 254820 96824
rect 255228 96772 255280 96824
rect 201868 96704 201920 96756
rect 206468 96704 206520 96756
rect 244280 96704 244332 96756
rect 245476 96704 245528 96756
rect 202696 96636 202748 96688
rect 208400 96636 208452 96688
rect 210424 96636 210476 96688
rect 216220 96636 216272 96688
rect 243084 96636 243136 96688
rect 246304 96636 246356 96688
rect 186964 96568 187016 96620
rect 231308 96568 231360 96620
rect 257068 96840 257120 96892
rect 257804 96840 257856 96892
rect 258816 96840 258868 96892
rect 259368 96840 259420 96892
rect 259644 96840 259696 96892
rect 260748 96840 260800 96892
rect 261668 96840 261720 96892
rect 262956 96840 263008 96892
rect 264244 96840 264296 96892
rect 264888 96840 264940 96892
rect 266636 96840 266688 96892
rect 267648 96840 267700 96892
rect 267832 96840 267884 96892
rect 268568 96840 268620 96892
rect 269580 96840 269632 96892
rect 270316 96840 270368 96892
rect 271972 96840 272024 96892
rect 273168 96840 273220 96892
rect 255412 96772 255464 96824
rect 256056 96772 256108 96824
rect 258264 96772 258316 96824
rect 259184 96772 259236 96824
rect 260196 96772 260248 96824
rect 260472 96772 260524 96824
rect 262404 96772 262456 96824
rect 263324 96772 263376 96824
rect 263784 96772 263836 96824
rect 264704 96772 264756 96824
rect 265624 96772 265676 96824
rect 266176 96772 266228 96824
rect 266452 96772 266504 96824
rect 267188 96772 267240 96824
rect 268384 96772 268436 96824
rect 268936 96772 268988 96824
rect 269396 96772 269448 96824
rect 270040 96772 270092 96824
rect 272156 96772 272208 96824
rect 273076 96772 273128 96824
rect 260012 96704 260064 96756
rect 260564 96704 260616 96756
rect 261392 96704 261444 96756
rect 262036 96704 262088 96756
rect 262220 96704 262272 96756
rect 263416 96704 263468 96756
rect 264980 96704 265032 96756
rect 266084 96704 266136 96756
rect 269212 96704 269264 96756
rect 270132 96704 270184 96756
rect 271880 96704 271932 96756
rect 274088 96772 274140 96824
rect 274364 96772 274416 96824
rect 277308 96840 277360 96892
rect 278136 96840 278188 96892
rect 278320 96840 278372 96892
rect 278504 96840 278556 96892
rect 279332 96840 279384 96892
rect 279976 96840 280028 96892
rect 280528 96840 280580 96892
rect 281172 96840 281224 96892
rect 281724 96840 281776 96892
rect 282644 96840 282696 96892
rect 283748 96840 283800 96892
rect 284116 96840 284168 96892
rect 284300 96840 284352 96892
rect 285496 96840 285548 96892
rect 285956 96840 286008 96892
rect 286692 96840 286744 96892
rect 273352 96704 273404 96756
rect 274640 96704 274692 96756
rect 275560 96704 275612 96756
rect 275836 96704 275888 96756
rect 276204 96704 276256 96756
rect 277308 96704 277360 96756
rect 260840 96636 260892 96688
rect 261944 96636 261996 96688
rect 273628 96636 273680 96688
rect 161388 96500 161440 96552
rect 206928 96500 206980 96552
rect 183468 96432 183520 96484
rect 230756 96432 230808 96484
rect 274824 96636 274876 96688
rect 276388 96636 276440 96688
rect 277216 96636 277268 96688
rect 277952 96772 278004 96824
rect 278688 96772 278740 96824
rect 278780 96772 278832 96824
rect 279884 96772 279936 96824
rect 280344 96772 280396 96824
rect 281264 96772 281316 96824
rect 282368 96772 282420 96824
rect 282552 96772 282604 96824
rect 283564 96772 283616 96824
rect 284024 96772 284076 96824
rect 286508 96772 286560 96824
rect 286784 96772 286836 96824
rect 277584 96704 277636 96756
rect 278596 96704 278648 96756
rect 279516 96704 279568 96756
rect 307024 96840 307076 96892
rect 287152 96772 287204 96824
rect 287796 96772 287848 96824
rect 289176 96772 289228 96824
rect 289728 96772 289780 96824
rect 290740 96772 290792 96824
rect 290924 96772 290976 96824
rect 291292 96772 291344 96824
rect 291936 96772 291988 96824
rect 292212 96772 292264 96824
rect 292488 96772 292540 96824
rect 294420 96772 294472 96824
rect 295248 96772 295300 96824
rect 295524 96772 295576 96824
rect 296444 96772 296496 96824
rect 296720 96772 296772 96824
rect 298100 96772 298152 96824
rect 298192 96772 298244 96824
rect 304356 96772 304408 96824
rect 287704 96704 287756 96756
rect 288072 96704 288124 96756
rect 288532 96704 288584 96756
rect 289544 96704 289596 96756
rect 291476 96704 291528 96756
rect 292120 96704 292172 96756
rect 294512 96704 294564 96756
rect 294972 96704 295024 96756
rect 296076 96704 296128 96756
rect 296352 96704 296404 96756
rect 296996 96704 297048 96756
rect 297824 96704 297876 96756
rect 298008 96704 298060 96756
rect 304264 96704 304316 96756
rect 282736 96636 282788 96688
rect 283104 96636 283156 96688
rect 283840 96636 283892 96688
rect 287336 96636 287388 96688
rect 287888 96636 287940 96688
rect 291844 96636 291896 96688
rect 292304 96636 292356 96688
rect 294144 96636 294196 96688
rect 294788 96636 294840 96688
rect 294880 96636 294932 96688
rect 295156 96636 295208 96688
rect 295708 96636 295760 96688
rect 296168 96636 296220 96688
rect 297272 96636 297324 96688
rect 297916 96636 297968 96688
rect 274364 96500 274416 96552
rect 275836 96500 275888 96552
rect 324964 96568 325016 96620
rect 285588 96500 285640 96552
rect 461584 96500 461636 96552
rect 283748 96432 283800 96484
rect 468484 96432 468536 96484
rect 179328 96364 179380 96416
rect 230112 96364 230164 96416
rect 285036 96364 285088 96416
rect 285404 96364 285456 96416
rect 176568 96296 176620 96348
rect 227720 96296 227772 96348
rect 282828 96296 282880 96348
rect 472624 96364 472676 96416
rect 173164 96228 173216 96280
rect 228916 96228 228968 96280
rect 282092 96228 282144 96280
rect 475384 96296 475436 96348
rect 285864 96228 285916 96280
rect 479524 96228 479576 96280
rect 169668 96160 169720 96212
rect 228364 96160 228416 96212
rect 281540 96160 281592 96212
rect 483020 96160 483072 96212
rect 155224 96092 155276 96144
rect 225972 96092 226024 96144
rect 283380 96092 283432 96144
rect 494060 96092 494112 96144
rect 133788 96024 133840 96076
rect 215300 96024 215352 96076
rect 284576 96024 284628 96076
rect 500960 96024 501012 96076
rect 70308 95956 70360 96008
rect 211620 95956 211672 96008
rect 280988 95956 281040 96008
rect 17868 95888 17920 95940
rect 202880 95888 202932 95940
rect 202972 95888 203024 95940
rect 203708 95888 203760 95940
rect 247684 95888 247736 95940
rect 282184 95888 282236 95940
rect 285772 95956 285824 96008
rect 507860 95956 507912 96008
rect 285864 95888 285916 95940
rect 297364 95888 297416 95940
rect 518900 95888 518952 95940
rect 165528 95820 165580 95872
rect 208124 95820 208176 95872
rect 253020 95820 253072 95872
rect 312544 95820 312596 95872
rect 191104 95752 191156 95804
rect 231952 95752 232004 95804
rect 252468 95752 252520 95804
rect 309140 95752 309192 95804
rect 197268 95684 197320 95736
rect 233148 95684 233200 95736
rect 242900 95684 242952 95736
rect 250444 95684 250496 95736
rect 251088 95684 251140 95736
rect 302240 95684 302292 95736
rect 200028 95616 200080 95668
rect 233884 95616 233936 95668
rect 256700 95616 256752 95668
rect 306380 95616 306432 95668
rect 194508 95548 194560 95600
rect 218060 95548 218112 95600
rect 249892 95548 249944 95600
rect 298192 95548 298244 95600
rect 262864 95480 262916 95532
rect 299480 95480 299532 95532
rect 287520 95412 287572 95464
rect 297364 95412 297416 95464
rect 233148 95344 233200 95396
rect 239128 95344 239180 95396
rect 234436 95276 234488 95328
rect 239956 95276 240008 95328
rect 228640 95208 228692 95260
rect 233976 95208 234028 95260
rect 162768 95140 162820 95192
rect 227352 95140 227404 95192
rect 286968 95140 287020 95192
rect 454684 95140 454736 95192
rect 158628 95072 158680 95124
rect 226524 95072 226576 95124
rect 279700 95072 279752 95124
rect 464344 95072 464396 95124
rect 144828 95004 144880 95056
rect 212540 95004 212592 95056
rect 292396 95004 292448 95056
rect 485044 95004 485096 95056
rect 147588 94936 147640 94988
rect 224776 94936 224828 94988
rect 291108 94936 291160 94988
rect 489184 94936 489236 94988
rect 137284 94868 137336 94920
rect 223028 94868 223080 94920
rect 289636 94868 289688 94920
rect 502984 94868 503036 94920
rect 128268 94800 128320 94852
rect 221372 94800 221424 94852
rect 286324 94800 286376 94852
rect 512000 94800 512052 94852
rect 78588 94732 78640 94784
rect 213092 94732 213144 94784
rect 288164 94732 288216 94784
rect 520924 94732 520976 94784
rect 64788 94664 64840 94716
rect 210792 94664 210844 94716
rect 229744 94664 229796 94716
rect 237564 94664 237616 94716
rect 288716 94664 288768 94716
rect 525800 94664 525852 94716
rect 37096 94596 37148 94648
rect 206284 94596 206336 94648
rect 244924 94596 244976 94648
rect 262864 94596 262916 94648
rect 290556 94596 290608 94648
rect 536840 94596 536892 94648
rect 33784 94528 33836 94580
rect 205272 94528 205324 94580
rect 208584 94528 208636 94580
rect 209504 94528 209556 94580
rect 210148 94528 210200 94580
rect 210608 94528 210660 94580
rect 212908 94528 212960 94580
rect 213552 94528 213604 94580
rect 214104 94528 214156 94580
rect 214748 94528 214800 94580
rect 233608 94528 233660 94580
rect 234252 94528 234304 94580
rect 248052 94528 248104 94580
rect 285680 94528 285732 94580
rect 291752 94528 291804 94580
rect 543740 94528 543792 94580
rect 25504 94460 25556 94512
rect 203616 94460 203668 94512
rect 209964 94460 210016 94512
rect 210884 94460 210936 94512
rect 224868 94460 224920 94512
rect 231860 94460 231912 94512
rect 249708 94460 249760 94512
rect 293224 94460 293276 94512
rect 293408 94460 293460 94512
rect 293776 94460 293828 94512
rect 295340 94460 295392 94512
rect 558184 94460 558236 94512
rect 166908 94392 166960 94444
rect 227996 94392 228048 94444
rect 230848 94392 230900 94444
rect 231676 94392 231728 94444
rect 259828 94392 259880 94444
rect 353944 94392 353996 94444
rect 157248 94324 157300 94376
rect 216680 94324 216732 94376
rect 231124 94324 231176 94376
rect 236920 94324 236972 94376
rect 255872 94324 255924 94376
rect 331220 94324 331272 94376
rect 174544 94256 174596 94308
rect 229192 94256 229244 94308
rect 253756 94256 253808 94308
rect 316040 94256 316092 94308
rect 177948 94188 178000 94240
rect 229652 94188 229704 94240
rect 252836 94188 252888 94240
rect 313280 94188 313332 94240
rect 184848 94120 184900 94172
rect 230756 94120 230808 94172
rect 262772 94120 262824 94172
rect 320180 94120 320232 94172
rect 198648 94052 198700 94104
rect 233240 94052 233292 94104
rect 292672 94052 292724 94104
rect 293684 94052 293736 94104
rect 160008 93780 160060 93832
rect 226800 93780 226852 93832
rect 261852 93780 261904 93832
rect 360844 93780 360896 93832
rect 155868 93712 155920 93764
rect 226064 93712 226116 93764
rect 262128 93712 262180 93764
rect 364984 93712 365036 93764
rect 148968 93644 149020 93696
rect 218796 93644 218848 93696
rect 263324 93644 263376 93696
rect 367744 93644 367796 93696
rect 153108 93576 153160 93628
rect 225420 93576 225472 93628
rect 264796 93576 264848 93628
rect 374644 93576 374696 93628
rect 144736 93508 144788 93560
rect 224040 93508 224092 93560
rect 270408 93508 270460 93560
rect 416780 93508 416832 93560
rect 142068 93440 142120 93492
rect 223672 93440 223724 93492
rect 273168 93440 273220 93492
rect 421564 93440 421616 93492
rect 131028 93372 131080 93424
rect 221464 93372 221516 93424
rect 275928 93372 275980 93424
rect 448520 93372 448572 93424
rect 84108 93304 84160 93356
rect 213828 93304 213880 93356
rect 293500 93304 293552 93356
rect 554044 93304 554096 93356
rect 73068 93236 73120 93288
rect 212080 93236 212132 93288
rect 294696 93236 294748 93288
rect 561680 93236 561732 93288
rect 68284 93168 68336 93220
rect 210056 93168 210108 93220
rect 243636 93168 243688 93220
rect 257344 93168 257396 93220
rect 295984 93168 296036 93220
rect 568580 93168 568632 93220
rect 14464 93100 14516 93152
rect 201500 93100 201552 93152
rect 246856 93100 246908 93152
rect 261484 93100 261536 93152
rect 296536 93100 296588 93152
rect 572720 93100 572772 93152
rect 170404 93032 170456 93084
rect 228456 93032 228508 93084
rect 257988 93032 258040 93084
rect 340880 93032 340932 93084
rect 180708 92964 180760 93016
rect 230204 92964 230256 93016
rect 257804 92964 257856 93016
rect 338120 92964 338172 93016
rect 188344 92896 188396 92948
rect 231400 92896 231452 92948
rect 256516 92896 256568 92948
rect 333980 92896 334032 92948
rect 229836 92556 229888 92608
rect 236552 92556 236604 92608
rect 231216 92488 231268 92540
rect 234620 92488 234672 92540
rect 177856 92420 177908 92472
rect 229928 92420 229980 92472
rect 264888 92420 264940 92472
rect 378784 92420 378836 92472
rect 175188 92352 175240 92404
rect 229376 92352 229428 92404
rect 264612 92352 264664 92404
rect 382924 92352 382976 92404
rect 169024 92284 169076 92336
rect 228180 92284 228232 92336
rect 267004 92284 267056 92336
rect 387800 92284 387852 92336
rect 164148 92216 164200 92268
rect 227444 92216 227496 92268
rect 266268 92216 266320 92268
rect 389824 92216 389876 92268
rect 128176 92148 128228 92200
rect 221556 92148 221608 92200
rect 272892 92148 272944 92200
rect 430580 92148 430632 92200
rect 104164 92080 104216 92132
rect 217048 92080 217100 92132
rect 272984 92080 273036 92132
rect 432604 92080 432656 92132
rect 79968 92012 80020 92064
rect 213276 92012 213328 92064
rect 277308 92012 277360 92064
rect 446404 92012 446456 92064
rect 77208 91944 77260 91996
rect 212816 91944 212868 91996
rect 277032 91944 277084 91996
rect 453304 91944 453356 91996
rect 54484 91876 54536 91928
rect 208492 91876 208544 91928
rect 278688 91876 278740 91928
rect 460204 91876 460256 91928
rect 45468 91808 45520 91860
rect 207480 91808 207532 91860
rect 246948 91808 247000 91860
rect 264244 91808 264296 91860
rect 279884 91808 279936 91860
rect 465724 91808 465776 91860
rect 23388 91740 23440 91792
rect 202972 91740 203024 91792
rect 230388 91740 230440 91792
rect 239404 91740 239456 91792
rect 244004 91740 244056 91792
rect 262220 91740 262272 91792
rect 287796 91740 287848 91792
rect 515404 91740 515456 91792
rect 182088 91672 182140 91724
rect 230664 91672 230716 91724
rect 233424 91672 233476 91724
rect 234068 91672 234120 91724
rect 260748 91672 260800 91724
rect 353300 91672 353352 91724
rect 187056 91604 187108 91656
rect 231032 91604 231084 91656
rect 256056 91604 256108 91656
rect 328460 91604 328512 91656
rect 232228 90992 232280 91044
rect 232596 90992 232648 91044
rect 274548 90992 274600 91044
rect 407764 90992 407816 91044
rect 153016 90924 153068 90976
rect 225696 90924 225748 90976
rect 269028 90924 269080 90976
rect 403624 90924 403676 90976
rect 146208 90856 146260 90908
rect 224500 90856 224552 90908
rect 289268 90856 289320 90908
rect 471244 90856 471296 90908
rect 112444 90788 112496 90840
rect 219072 90788 219124 90840
rect 278412 90788 278464 90840
rect 465172 90788 465224 90840
rect 108948 90720 109000 90772
rect 218888 90720 218940 90772
rect 282644 90720 282696 90772
rect 476764 90720 476816 90772
rect 105544 90652 105596 90704
rect 217508 90652 217560 90704
rect 282552 90652 282604 90704
rect 486424 90652 486476 90704
rect 90364 90584 90416 90636
rect 214932 90584 214984 90636
rect 284024 90584 284076 90636
rect 493324 90584 493376 90636
rect 75184 90516 75236 90568
rect 211344 90516 211396 90568
rect 283932 90516 283984 90568
rect 497464 90516 497516 90568
rect 65524 90448 65576 90500
rect 209320 90448 209372 90500
rect 285128 90448 285180 90500
rect 500224 90448 500276 90500
rect 53104 90380 53156 90432
rect 208032 90380 208084 90432
rect 286692 90380 286744 90432
rect 504364 90380 504416 90432
rect 41328 90312 41380 90364
rect 206744 90312 206796 90364
rect 217324 90312 217376 90364
rect 234344 90312 234396 90364
rect 244096 90312 244148 90364
rect 255964 90312 256016 90364
rect 291936 90312 291988 90364
rect 540244 90312 540296 90364
rect 263416 90244 263468 90296
rect 356704 90244 356756 90296
rect 257896 90176 257948 90228
rect 339500 90176 339552 90228
rect 256332 90108 256384 90160
rect 335360 90108 335412 90160
rect 253572 90040 253624 90092
rect 317420 90040 317472 90092
rect 259000 89632 259052 89684
rect 346400 89632 346452 89684
rect 265992 89564 266044 89616
rect 385684 89564 385736 89616
rect 124128 89496 124180 89548
rect 221280 89496 221332 89548
rect 271696 89496 271748 89548
rect 410524 89496 410576 89548
rect 116584 89428 116636 89480
rect 218520 89428 218572 89480
rect 275652 89428 275704 89480
rect 442264 89428 442316 89480
rect 103428 89360 103480 89412
rect 216864 89360 216916 89412
rect 285312 89360 285364 89412
rect 506480 89360 506532 89412
rect 80704 89292 80756 89344
rect 211712 89292 211764 89344
rect 286784 89292 286836 89344
rect 511264 89292 511316 89344
rect 79324 89224 79376 89276
rect 213000 89224 213052 89276
rect 288072 89224 288124 89276
rect 518164 89224 518216 89276
rect 70216 89156 70268 89208
rect 211528 89156 211580 89208
rect 288256 89156 288308 89208
rect 522304 89156 522356 89208
rect 47584 89088 47636 89140
rect 204720 89088 204772 89140
rect 289452 89088 289504 89140
rect 529204 89088 529256 89140
rect 35164 89020 35216 89072
rect 203156 89020 203208 89072
rect 290924 89020 290976 89072
rect 538220 89020 538272 89072
rect 21364 88952 21416 89004
rect 201776 88952 201828 89004
rect 248144 88952 248196 89004
rect 287060 88952 287112 89004
rect 296352 88952 296404 89004
rect 569960 88952 570012 89004
rect 257712 88884 257764 88936
rect 342260 88884 342312 88936
rect 256424 88816 256476 88868
rect 331864 88816 331916 88868
rect 253664 88748 253716 88800
rect 311256 88748 311308 88800
rect 261944 88272 261996 88324
rect 360200 88272 360252 88324
rect 262036 88204 262088 88256
rect 364340 88204 364392 88256
rect 263508 88136 263560 88188
rect 374092 88136 374144 88188
rect 264704 88068 264756 88120
rect 378140 88068 378192 88120
rect 267188 88000 267240 88052
rect 392584 88000 392636 88052
rect 111064 87932 111116 87984
rect 218336 87932 218388 87984
rect 273076 87932 273128 87984
rect 427820 87932 427872 87984
rect 88984 87864 89036 87916
rect 208952 87864 209004 87916
rect 274180 87864 274232 87916
rect 438860 87864 438912 87916
rect 87604 87796 87656 87848
rect 208584 87796 208636 87848
rect 293684 87796 293736 87848
rect 536104 87796 536156 87848
rect 86224 87728 86276 87780
rect 212908 87728 212960 87780
rect 292304 87728 292356 87780
rect 543004 87728 543056 87780
rect 44088 87660 44140 87712
rect 203524 87660 203576 87712
rect 292212 87660 292264 87712
rect 547972 87660 548024 87712
rect 15844 87592 15896 87644
rect 202328 87592 202380 87644
rect 296444 87592 296496 87644
rect 565820 87592 565872 87644
rect 260472 87524 260524 87576
rect 357440 87524 357492 87576
rect 311164 86912 311216 86964
rect 580172 86912 580224 86964
rect 261760 86844 261812 86896
rect 367100 86844 367152 86896
rect 270040 86776 270092 86828
rect 381544 86776 381596 86828
rect 264428 86708 264480 86760
rect 382372 86708 382424 86760
rect 267280 86640 267332 86692
rect 395344 86640 395396 86692
rect 272800 86572 272852 86624
rect 406384 86572 406436 86624
rect 274272 86504 274324 86556
rect 441620 86504 441672 86556
rect 122104 86436 122156 86488
rect 217416 86436 217468 86488
rect 275744 86436 275796 86488
rect 448612 86436 448664 86488
rect 33048 86368 33100 86420
rect 199384 86368 199436 86420
rect 279976 86368 280028 86420
rect 470600 86368 470652 86420
rect 28264 86300 28316 86352
rect 201592 86300 201644 86352
rect 284116 86300 284168 86352
rect 496820 86300 496872 86352
rect 5448 86232 5500 86284
rect 195336 86232 195388 86284
rect 290464 86232 290516 86284
rect 535460 86232 535512 86284
rect 256148 86164 256200 86216
rect 329840 86164 329892 86216
rect 3148 85484 3200 85536
rect 151084 85484 151136 85536
rect 253388 85416 253440 85468
rect 318064 85416 318116 85468
rect 263048 85348 263100 85400
rect 340972 85348 341024 85400
rect 259092 85280 259144 85332
rect 342904 85280 342956 85332
rect 271328 85212 271380 85264
rect 375380 85212 375432 85264
rect 279792 85144 279844 85196
rect 472716 85144 472768 85196
rect 281908 85076 281960 85128
rect 482284 85076 482336 85128
rect 283840 85008 283892 85060
rect 492680 85008 492732 85060
rect 285496 84940 285548 84992
rect 499580 84940 499632 84992
rect 289544 84872 289596 84924
rect 524420 84872 524472 84924
rect 107568 84804 107620 84856
rect 196624 84804 196676 84856
rect 293776 84804 293828 84856
rect 553400 84804 553452 84856
rect 276664 83852 276716 83904
rect 357532 83852 357584 83904
rect 262956 83784 263008 83836
rect 365812 83784 365864 83836
rect 274364 83716 274416 83768
rect 418804 83716 418856 83768
rect 286508 83648 286560 83700
rect 510620 83648 510672 83700
rect 287888 83580 287940 83632
rect 517520 83580 517572 83632
rect 290832 83512 290884 83564
rect 539692 83512 539744 83564
rect 246672 83444 246724 83496
rect 273904 83444 273956 83496
rect 293592 83444 293644 83496
rect 556252 83444 556304 83496
rect 298836 82424 298888 82476
rect 400220 82424 400272 82476
rect 264520 82356 264572 82408
rect 377404 82356 377456 82408
rect 275836 82288 275888 82340
rect 396724 82288 396776 82340
rect 271788 82220 271840 82272
rect 393964 82220 394016 82272
rect 296168 82152 296220 82204
rect 565084 82152 565136 82204
rect 248236 82084 248288 82136
rect 275284 82084 275336 82136
rect 278504 82084 278556 82136
rect 295984 82084 296036 82136
rect 304356 82084 304408 82136
rect 582564 82084 582616 82136
rect 275560 80792 275612 80844
rect 399484 80792 399536 80844
rect 274456 80724 274508 80776
rect 411904 80724 411956 80776
rect 248052 80656 248104 80708
rect 284300 80656 284352 80708
rect 298744 80656 298796 80708
rect 575480 80656 575532 80708
rect 316684 73108 316736 73160
rect 579988 73108 580040 73160
rect 253480 72428 253532 72480
rect 316132 72428 316184 72480
rect 3424 71680 3476 71732
rect 157984 71680 158036 71732
rect 530584 60664 530636 60716
rect 580172 60664 580224 60716
rect 289176 59984 289228 60036
rect 530676 59984 530728 60036
rect 3056 59304 3108 59356
rect 32404 59304 32456 59356
rect 68928 47540 68980 47592
rect 198004 47540 198056 47592
rect 3424 45500 3476 45552
rect 148324 45500 148376 45552
rect 3148 33056 3200 33108
rect 156604 33056 156656 33108
rect 313924 33056 313976 33108
rect 580172 33056 580224 33108
rect 286600 26868 286652 26920
rect 514852 26868 514904 26920
rect 285036 24080 285088 24132
rect 506572 24080 506624 24132
rect 296260 22720 296312 22772
rect 571340 22720 571392 22772
rect 292028 21360 292080 21412
rect 546500 21360 546552 21412
rect 3424 20612 3476 20664
rect 43444 20612 43496 20664
rect 525064 20612 525116 20664
rect 580172 20612 580224 20664
rect 282460 19932 282512 19984
rect 490012 19932 490064 19984
rect 188988 18572 189040 18624
rect 230848 18572 230900 18624
rect 287980 18572 288032 18624
rect 521660 18572 521712 18624
rect 250812 16056 250864 16108
rect 298100 16056 298152 16108
rect 250904 15988 250956 16040
rect 301504 15988 301556 16040
rect 252100 15920 252152 15972
rect 307760 15920 307812 15972
rect 106188 15852 106240 15904
rect 217140 15852 217192 15904
rect 240048 15852 240100 15904
rect 253480 15852 253532 15904
rect 254860 15852 254912 15904
rect 322940 15852 322992 15904
rect 323584 15852 323636 15904
rect 404360 15852 404412 15904
rect 294972 14628 295024 14680
rect 560392 14628 560444 14680
rect 294880 14560 294932 14612
rect 564440 14560 564492 14612
rect 297824 14492 297876 14544
rect 575112 14492 575164 14544
rect 161204 14424 161256 14476
rect 226616 14424 226668 14476
rect 258724 14424 258776 14476
rect 281540 14424 281592 14476
rect 297732 14424 297784 14476
rect 578608 14424 578660 14476
rect 256240 13472 256292 13524
rect 333888 13472 333940 13524
rect 277216 13404 277268 13456
rect 453212 13404 453264 13456
rect 277124 13336 277176 13388
rect 456892 13336 456944 13388
rect 278596 13268 278648 13320
rect 459928 13268 459980 13320
rect 278320 13200 278372 13252
rect 463976 13200 464028 13252
rect 281172 13132 281224 13184
rect 478144 13132 478196 13184
rect 170772 13064 170824 13116
rect 228088 13064 228140 13116
rect 246764 13064 246816 13116
rect 267004 13064 267056 13116
rect 281080 13064 281132 13116
rect 482192 13064 482244 13116
rect 266084 12248 266136 12300
rect 385592 12248 385644 12300
rect 266176 12180 266228 12232
rect 389456 12180 389508 12232
rect 265900 12112 265952 12164
rect 392584 12112 392636 12164
rect 267372 12044 267424 12096
rect 396080 12044 396132 12096
rect 267464 11976 267516 12028
rect 398840 11976 398892 12028
rect 268660 11908 268712 11960
rect 403532 11908 403584 11960
rect 268752 11840 268804 11892
rect 407212 11840 407264 11892
rect 245200 11772 245252 11824
rect 256056 11772 256108 11824
rect 270132 11772 270184 11824
rect 410432 11772 410484 11824
rect 111708 11704 111760 11756
rect 119344 11704 119396 11756
rect 119896 11704 119948 11756
rect 219900 11704 219952 11756
rect 243912 11704 243964 11756
rect 256148 11704 256200 11756
rect 270224 11704 270276 11756
rect 414296 11704 414348 11756
rect 357532 11636 357584 11688
rect 358728 11636 358780 11688
rect 250996 10888 251048 10940
rect 299572 10888 299624 10940
rect 252192 10820 252244 10872
rect 303896 10820 303948 10872
rect 252284 10752 252336 10804
rect 307944 10752 307996 10804
rect 252376 10684 252428 10736
rect 311164 10684 311216 10736
rect 117228 10616 117280 10668
rect 220268 10616 220320 10668
rect 255044 10616 255096 10668
rect 322112 10616 322164 10668
rect 99288 10548 99340 10600
rect 215484 10548 215536 10600
rect 254952 10548 255004 10600
rect 324320 10548 324372 10600
rect 95148 10480 95200 10532
rect 216036 10480 216088 10532
rect 295156 10480 295208 10532
rect 559288 10480 559340 10532
rect 92388 10412 92440 10464
rect 215668 10412 215720 10464
rect 295064 10412 295116 10464
rect 563244 10412 563296 10464
rect 87972 10344 88024 10396
rect 214104 10344 214156 10396
rect 298008 10344 298060 10396
rect 573456 10344 573508 10396
rect 85488 10276 85540 10328
rect 214196 10276 214248 10328
rect 297916 10276 297968 10328
rect 576952 10276 577004 10328
rect 122288 9460 122340 9512
rect 219716 9460 219768 9512
rect 118792 9392 118844 9444
rect 219532 9392 219584 9444
rect 115296 9324 115348 9376
rect 220452 9324 220504 9376
rect 97448 9256 97500 9308
rect 215760 9256 215812 9308
rect 93952 9188 94004 9240
rect 215852 9188 215904 9240
rect 90456 9120 90508 9172
rect 214472 9120 214524 9172
rect 86868 9052 86920 9104
rect 214288 9052 214340 9104
rect 300124 9052 300176 9104
rect 362316 9052 362368 9104
rect 33600 8984 33652 9036
rect 205640 8984 205692 9036
rect 281264 8984 281316 9036
rect 476948 8984 477000 9036
rect 30104 8916 30156 8968
rect 204996 8916 205048 8968
rect 220452 8916 220504 8968
rect 231308 8916 231360 8968
rect 253204 8916 253256 8968
rect 280712 8916 280764 8968
rect 281356 8916 281408 8968
rect 481732 8916 481784 8968
rect 260104 8236 260156 8288
rect 264152 8236 264204 8288
rect 202696 8100 202748 8152
rect 233424 8100 233476 8152
rect 199108 8032 199160 8084
rect 233792 8032 233844 8084
rect 267648 8032 267700 8084
rect 395252 8032 395304 8084
rect 75000 7896 75052 7948
rect 142804 7964 142856 8016
rect 195612 7964 195664 8016
rect 232688 7964 232740 8016
rect 267556 7964 267608 8016
rect 398932 7964 398984 8016
rect 142436 7896 142488 7948
rect 223948 7896 224000 7948
rect 268568 7896 268620 7948
rect 402520 7896 402572 7948
rect 138848 7760 138900 7812
rect 222476 7828 222528 7880
rect 268936 7828 268988 7880
rect 406016 7828 406068 7880
rect 146944 7760 146996 7812
rect 222752 7760 222804 7812
rect 268844 7760 268896 7812
rect 409604 7760 409656 7812
rect 131764 7692 131816 7744
rect 222936 7692 222988 7744
rect 270316 7692 270368 7744
rect 413100 7692 413152 7744
rect 50160 7624 50212 7676
rect 192484 7624 192536 7676
rect 192576 7624 192628 7676
rect 232044 7624 232096 7676
rect 269948 7624 270000 7676
rect 416688 7624 416740 7676
rect 26516 7556 26568 7608
rect 204352 7556 204404 7608
rect 209780 7556 209832 7608
rect 235080 7556 235132 7608
rect 249984 7556 250036 7608
rect 258448 7556 258500 7608
rect 274088 7556 274140 7608
rect 441528 7556 441580 7608
rect 448612 7556 448664 7608
rect 449808 7556 449860 7608
rect 135260 7488 135312 7540
rect 146944 7488 146996 7540
rect 3424 6808 3476 6860
rect 26884 6808 26936 6860
rect 249340 6672 249392 6724
rect 287796 6672 287848 6724
rect 194416 6604 194468 6656
rect 232228 6604 232280 6656
rect 255136 6604 255188 6656
rect 324412 6604 324464 6656
rect 190828 6536 190880 6588
rect 232412 6536 232464 6588
rect 254768 6536 254820 6588
rect 328000 6536 328052 6588
rect 134156 6468 134208 6520
rect 85672 6400 85724 6452
rect 134524 6400 134576 6452
rect 137652 6468 137704 6520
rect 222292 6468 222344 6520
rect 259184 6468 259236 6520
rect 345756 6468 345808 6520
rect 222660 6400 222712 6452
rect 260288 6400 260340 6452
rect 352840 6536 352892 6588
rect 65616 6332 65668 6384
rect 209964 6332 210016 6384
rect 260564 6332 260616 6384
rect 356336 6468 356388 6520
rect 352564 6400 352616 6452
rect 418988 6400 419040 6452
rect 62028 6264 62080 6316
rect 210700 6264 210752 6316
rect 215668 6264 215720 6316
rect 236276 6264 236328 6316
rect 260380 6264 260432 6316
rect 359924 6332 359976 6384
rect 359464 6264 359516 6316
rect 426164 6332 426216 6384
rect 425704 6264 425756 6316
rect 447416 6264 447468 6316
rect 447784 6264 447836 6316
rect 475752 6264 475804 6316
rect 38384 6196 38436 6248
rect 195244 6196 195296 6248
rect 212172 6196 212224 6248
rect 235632 6196 235684 6248
rect 250720 6196 250772 6248
rect 297272 6196 297324 6248
rect 307024 6196 307076 6248
rect 472256 6196 472308 6248
rect 4068 6128 4120 6180
rect 200580 6128 200632 6180
rect 208584 6128 208636 6180
rect 234988 6128 235040 6180
rect 249248 6128 249300 6180
rect 291384 6128 291436 6180
rect 292120 6128 292172 6180
rect 543188 6128 543240 6180
rect 234620 5516 234672 5568
rect 239036 5516 239088 5568
rect 24216 5176 24268 5228
rect 98644 5176 98696 5228
rect 99840 5176 99892 5228
rect 124864 5244 124916 5296
rect 245384 5176 245436 5228
rect 265348 5176 265400 5228
rect 370504 5176 370556 5228
rect 433248 5176 433300 5228
rect 35992 5108 36044 5160
rect 58624 5108 58676 5160
rect 58716 5108 58768 5160
rect 209872 5108 209924 5160
rect 249156 5108 249208 5160
rect 290188 5108 290240 5160
rect 363604 5108 363656 5160
rect 429660 5108 429712 5160
rect 54944 5040 54996 5092
rect 208952 5040 209004 5092
rect 221556 5040 221608 5092
rect 236460 5040 236512 5092
rect 249616 5040 249668 5092
rect 293684 5040 293736 5092
rect 302884 5040 302936 5092
rect 372896 5040 372948 5092
rect 429844 5040 429896 5092
rect 454500 5040 454552 5092
rect 47860 4972 47912 5024
rect 207296 4972 207348 5024
rect 218060 4972 218112 5024
rect 236644 4972 236696 5024
rect 245292 4972 245344 5024
rect 268844 4972 268896 5024
rect 271236 4972 271288 5024
rect 415492 4972 415544 5024
rect 450544 4972 450596 5024
rect 582196 4972 582248 5024
rect 2872 4904 2924 4956
rect 200396 4904 200448 4956
rect 214472 4904 214524 4956
rect 236184 4904 236236 4956
rect 246488 4904 246540 4956
rect 276020 4904 276072 4956
rect 285220 4904 285272 4956
rect 504180 4904 504232 4956
rect 1676 4836 1728 4888
rect 200304 4836 200356 4888
rect 210976 4836 211028 4888
rect 235540 4836 235592 4888
rect 249524 4836 249576 4888
rect 288992 4836 289044 4888
rect 289360 4836 289412 4888
rect 529020 4836 529072 4888
rect 572 4768 624 4820
rect 200120 4768 200172 4820
rect 207388 4768 207440 4820
rect 234804 4768 234856 4820
rect 249432 4768 249484 4820
rect 292580 4768 292632 4820
rect 294788 4768 294840 4820
rect 558552 4768 558604 4820
rect 60832 4088 60884 4140
rect 71044 4088 71096 4140
rect 73804 4088 73856 4140
rect 80704 4088 80756 4140
rect 82084 4088 82136 4140
rect 124680 4156 124732 4208
rect 126244 4156 126296 4208
rect 241244 4156 241296 4208
rect 242900 4156 242952 4208
rect 93124 4088 93176 4140
rect 146944 4088 146996 4140
rect 223580 4088 223632 4140
rect 228732 4088 228784 4140
rect 237656 4088 237708 4140
rect 257344 4088 257396 4140
rect 258264 4088 258316 4140
rect 353944 4088 353996 4140
rect 355232 4088 355284 4140
rect 410524 4088 410576 4140
rect 424968 4088 425020 4140
rect 453304 4088 453356 4140
rect 455696 4088 455748 4140
rect 460204 4088 460256 4140
rect 462780 4088 462832 4140
rect 479524 4088 479576 4140
rect 480536 4088 480588 4140
rect 518164 4088 518216 4140
rect 520740 4088 520792 4140
rect 565084 4088 565136 4140
rect 568028 4088 568080 4140
rect 34796 4020 34848 4072
rect 46204 4020 46256 4072
rect 57244 4020 57296 4072
rect 87604 4020 87656 4072
rect 101036 4020 101088 4072
rect 104164 4020 104216 4072
rect 19432 3952 19484 4004
rect 35164 3952 35216 4004
rect 56048 3952 56100 4004
rect 65524 3952 65576 4004
rect 71504 3952 71556 4004
rect 101404 3952 101456 4004
rect 103336 3952 103388 4004
rect 122104 4020 122156 4072
rect 129372 4020 129424 4072
rect 221096 4020 221148 4072
rect 117596 3952 117648 4004
rect 214564 3952 214616 4004
rect 223764 3952 223816 4004
rect 228364 3952 228416 4004
rect 28908 3884 28960 3936
rect 47584 3884 47636 3936
rect 53748 3884 53800 3936
rect 88984 3884 89036 3936
rect 92756 3884 92808 3936
rect 97264 3884 97316 3936
rect 112812 3884 112864 3936
rect 116584 3884 116636 3936
rect 121092 3884 121144 3936
rect 220084 3884 220136 3936
rect 226340 3884 226392 3936
rect 238208 4020 238260 4072
rect 256148 4020 256200 4072
rect 260656 4020 260708 4072
rect 406384 4020 406436 4072
rect 259276 3952 259328 4004
rect 266728 3952 266780 4004
rect 267004 3952 267056 4004
rect 271236 3952 271288 4004
rect 273904 3952 273956 4004
rect 278320 3952 278372 4004
rect 296076 3952 296128 4004
rect 298192 3952 298244 4004
rect 392676 3952 392728 4004
rect 394240 3952 394292 4004
rect 418804 4020 418856 4072
rect 436744 4020 436796 4072
rect 464344 4020 464396 4072
rect 473452 4020 473504 4072
rect 432052 3952 432104 4004
rect 436836 3952 436888 4004
rect 11152 3816 11204 3868
rect 28264 3816 28316 3868
rect 46664 3816 46716 3868
rect 94504 3816 94556 3868
rect 96252 3816 96304 3868
rect 210424 3816 210476 3868
rect 225144 3816 225196 3868
rect 237932 3884 237984 3936
rect 256056 3884 256108 3936
rect 267740 3884 267792 3936
rect 304264 3884 304316 3936
rect 351644 3884 351696 3936
rect 407764 3884 407816 3936
rect 435548 3884 435600 3936
rect 229928 3816 229980 3868
rect 238116 3816 238168 3868
rect 242808 3816 242860 3868
rect 251180 3816 251232 3868
rect 255964 3816 256016 3868
rect 259460 3816 259512 3868
rect 261484 3816 261536 3868
rect 277124 3816 277176 3868
rect 299572 3816 299624 3868
rect 300768 3816 300820 3868
rect 322204 3816 322256 3868
rect 383568 3816 383620 3868
rect 393964 3816 394016 3868
rect 422576 3816 422628 3868
rect 440884 3816 440936 3868
rect 445024 3816 445076 3868
rect 476764 3952 476816 4004
rect 485228 3952 485280 4004
rect 472624 3884 472676 3936
rect 491116 3884 491168 3936
rect 461584 3816 461636 3868
rect 468484 3816 468536 3868
rect 498200 3816 498252 3868
rect 503076 3816 503128 3868
rect 530124 3816 530176 3868
rect 20628 3748 20680 3800
rect 39304 3748 39356 3800
rect 45376 3748 45428 3800
rect 57152 3748 57204 3800
rect 63224 3748 63276 3800
rect 210148 3748 210200 3800
rect 219256 3748 219308 3800
rect 231124 3748 231176 3800
rect 252008 3748 252060 3800
rect 13544 3680 13596 3732
rect 36544 3680 36596 3732
rect 41880 3680 41932 3732
rect 50344 3680 50396 3732
rect 51356 3680 51408 3732
rect 208768 3680 208820 3732
rect 216864 3680 216916 3732
rect 229836 3680 229888 3732
rect 242624 3680 242676 3732
rect 252376 3680 252428 3732
rect 259368 3748 259420 3800
rect 349252 3748 349304 3800
rect 381544 3748 381596 3800
rect 411904 3748 411956 3800
rect 411996 3748 412048 3800
rect 440332 3748 440384 3800
rect 443644 3748 443696 3800
rect 305552 3680 305604 3732
rect 327724 3680 327776 3732
rect 390652 3680 390704 3732
rect 396724 3680 396776 3732
rect 443828 3680 443880 3732
rect 461676 3748 461728 3800
rect 505376 3748 505428 3800
rect 468668 3680 468720 3732
rect 475384 3680 475436 3732
rect 487620 3680 487672 3732
rect 489184 3680 489236 3732
rect 540796 3680 540848 3732
rect 9956 3612 10008 3664
rect 21364 3612 21416 3664
rect 25320 3612 25372 3664
rect 204260 3612 204312 3664
rect 213368 3612 213420 3664
rect 231216 3612 231268 3664
rect 238116 3612 238168 3664
rect 240968 3612 241020 3664
rect 246304 3612 246356 3664
rect 255872 3612 255924 3664
rect 7656 3544 7708 3596
rect 14740 3476 14792 3528
rect 15844 3476 15896 3528
rect 17040 3544 17092 3596
rect 17868 3544 17920 3596
rect 18236 3544 18288 3596
rect 19248 3544 19300 3596
rect 21824 3544 21876 3596
rect 25504 3544 25556 3596
rect 27712 3544 27764 3596
rect 29644 3544 29696 3596
rect 32404 3544 32456 3596
rect 33048 3544 33100 3596
rect 40684 3544 40736 3596
rect 41328 3544 41380 3596
rect 43076 3544 43128 3596
rect 44088 3544 44140 3596
rect 44272 3544 44324 3596
rect 45468 3544 45520 3596
rect 52552 3544 52604 3596
rect 54484 3544 54536 3596
rect 64328 3544 64380 3596
rect 64788 3544 64840 3596
rect 67916 3544 67968 3596
rect 68928 3544 68980 3596
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 72608 3544 72660 3596
rect 73068 3544 73120 3596
rect 76196 3544 76248 3596
rect 77208 3544 77260 3596
rect 77392 3544 77444 3596
rect 79324 3544 79376 3596
rect 83280 3544 83332 3596
rect 84108 3544 84160 3596
rect 84476 3544 84528 3596
rect 85488 3544 85540 3596
rect 89168 3544 89220 3596
rect 90364 3544 90416 3596
rect 91560 3544 91612 3596
rect 92388 3544 92440 3596
rect 98644 3544 98696 3596
rect 99288 3544 99340 3596
rect 102232 3544 102284 3596
rect 103428 3544 103480 3596
rect 105728 3544 105780 3596
rect 106188 3544 106240 3596
rect 106924 3544 106976 3596
rect 107568 3544 107620 3596
rect 108120 3544 108172 3596
rect 108948 3544 109000 3596
rect 109316 3544 109368 3596
rect 111064 3544 111116 3596
rect 111616 3544 111668 3596
rect 112444 3544 112496 3596
rect 114008 3544 114060 3596
rect 115204 3544 115256 3596
rect 116400 3544 116452 3596
rect 117228 3544 117280 3596
rect 123484 3544 123536 3596
rect 124128 3544 124180 3596
rect 125876 3544 125928 3596
rect 126888 3544 126940 3596
rect 126980 3544 127032 3596
rect 128268 3544 128320 3596
rect 130568 3544 130620 3596
rect 131028 3544 131080 3596
rect 132960 3544 133012 3596
rect 133788 3544 133840 3596
rect 136456 3544 136508 3596
rect 137284 3544 137336 3596
rect 140044 3544 140096 3596
rect 146944 3544 146996 3596
rect 147128 3544 147180 3596
rect 147588 3544 147640 3596
rect 148324 3544 148376 3596
rect 148968 3544 149020 3596
rect 149520 3544 149572 3596
rect 150348 3544 150400 3596
rect 151820 3544 151872 3596
rect 153108 3544 153160 3596
rect 154212 3544 154264 3596
rect 155224 3544 155276 3596
rect 155408 3544 155460 3596
rect 155868 3544 155920 3596
rect 156604 3544 156656 3596
rect 157248 3544 157300 3596
rect 157800 3544 157852 3596
rect 158628 3544 158680 3596
rect 158904 3544 158956 3596
rect 160008 3544 160060 3596
rect 160100 3544 160152 3596
rect 161204 3544 161256 3596
rect 163688 3544 163740 3596
rect 164148 3544 164200 3596
rect 164884 3544 164936 3596
rect 165528 3544 165580 3596
rect 166080 3544 166132 3596
rect 166908 3544 166960 3596
rect 167184 3544 167236 3596
rect 169024 3544 169076 3596
rect 171968 3544 172020 3596
rect 173164 3544 173216 3596
rect 174268 3544 174320 3596
rect 175188 3544 175240 3596
rect 175464 3544 175516 3596
rect 176568 3544 176620 3596
rect 176660 3544 176712 3596
rect 177948 3544 178000 3596
rect 180248 3544 180300 3596
rect 180708 3544 180760 3596
rect 181444 3544 181496 3596
rect 182088 3544 182140 3596
rect 182548 3544 182600 3596
rect 183468 3544 183520 3596
rect 183744 3544 183796 3596
rect 184848 3544 184900 3596
rect 186136 3544 186188 3596
rect 186964 3544 187016 3596
rect 187332 3544 187384 3596
rect 188344 3544 188396 3596
rect 188528 3544 188580 3596
rect 188988 3544 189040 3596
rect 189724 3544 189776 3596
rect 191104 3544 191156 3596
rect 192024 3544 192076 3596
rect 192576 3544 192628 3596
rect 193220 3544 193272 3596
rect 194508 3544 194560 3596
rect 196808 3544 196860 3596
rect 197268 3544 197320 3596
rect 197912 3544 197964 3596
rect 198648 3544 198700 3596
rect 201500 3544 201552 3596
rect 223764 3544 223816 3596
rect 200948 3476 201000 3528
rect 206192 3476 206244 3528
rect 235448 3544 235500 3596
rect 241428 3544 241480 3596
rect 244096 3544 244148 3596
rect 245476 3544 245528 3596
rect 262956 3612 263008 3664
rect 264244 3612 264296 3664
rect 261760 3544 261812 3596
rect 262220 3544 262272 3596
rect 262864 3544 262916 3596
rect 266544 3544 266596 3596
rect 266728 3612 266780 3664
rect 350448 3612 350500 3664
rect 356704 3612 356756 3664
rect 369400 3612 369452 3664
rect 395344 3612 395396 3664
rect 397736 3612 397788 3664
rect 399484 3612 399536 3664
rect 450912 3612 450964 3664
rect 454684 3612 454736 3664
rect 515956 3612 516008 3664
rect 273628 3544 273680 3596
rect 293224 3544 293276 3596
rect 294880 3544 294932 3596
rect 295984 3544 296036 3596
rect 465172 3544 465224 3596
rect 467104 3544 467156 3596
rect 469864 3544 469916 3596
rect 471244 3544 471296 3596
rect 527824 3612 527876 3664
rect 520924 3544 520976 3596
rect 523040 3544 523092 3596
rect 540244 3544 540296 3596
rect 541992 3544 542044 3596
rect 547144 3544 547196 3596
rect 552664 3544 552716 3596
rect 223948 3476 224000 3528
rect 224868 3476 224920 3528
rect 230388 3476 230440 3528
rect 231032 3476 231084 3528
rect 232228 3476 232280 3528
rect 233148 3476 233200 3528
rect 245108 3476 245160 3528
rect 270040 3476 270092 3528
rect 271144 3476 271196 3528
rect 274824 3476 274876 3528
rect 276940 3476 276992 3528
rect 449164 3476 449216 3528
rect 6460 3408 6512 3460
rect 200396 3408 200448 3460
rect 203892 3408 203944 3460
rect 233608 3408 233660 3460
rect 234436 3408 234488 3460
rect 237012 3408 237064 3460
rect 246580 3408 246632 3460
rect 272432 3408 272484 3460
rect 282184 3408 282236 3460
rect 283104 3408 283156 3460
rect 457444 3476 457496 3528
rect 534908 3476 534960 3528
rect 536104 3476 536156 3528
rect 550272 3476 550324 3528
rect 66720 3340 66772 3392
rect 75184 3340 75236 3392
rect 80888 3340 80940 3392
rect 86224 3340 86276 3392
rect 110512 3340 110564 3392
rect 111708 3340 111760 3392
rect 141240 3340 141292 3392
rect 142068 3340 142120 3392
rect 150624 3340 150676 3392
rect 225236 3340 225288 3392
rect 242716 3340 242768 3392
rect 59636 3272 59688 3324
rect 68284 3272 68336 3324
rect 169576 3272 169628 3324
rect 170404 3272 170456 3324
rect 205088 3272 205140 3324
rect 217324 3272 217376 3324
rect 242440 3272 242492 3324
rect 246396 3272 246448 3324
rect 280988 3340 281040 3392
rect 479340 3408 479392 3460
rect 486424 3408 486476 3460
rect 488816 3408 488868 3460
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 311256 3340 311308 3392
rect 312636 3340 312688 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 318156 3340 318208 3392
rect 319720 3340 319772 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 331864 3340 331916 3392
rect 332692 3340 332744 3392
rect 336004 3340 336056 3392
rect 337476 3340 337528 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 342996 3340 343048 3392
rect 344560 3340 344612 3392
rect 345664 3340 345716 3392
rect 348056 3340 348108 3392
rect 360844 3340 360896 3392
rect 363512 3340 363564 3392
rect 367836 3340 367888 3392
rect 370596 3340 370648 3392
rect 374644 3340 374696 3392
rect 377680 3340 377732 3392
rect 378784 3340 378836 3392
rect 381176 3340 381228 3392
rect 382924 3340 382976 3392
rect 384764 3340 384816 3392
rect 389824 3340 389876 3392
rect 391848 3340 391900 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 403624 3340 403676 3392
rect 408408 3340 408460 3392
rect 414664 3340 414716 3392
rect 421380 3340 421432 3392
rect 421564 3340 421616 3392
rect 427268 3340 427320 3392
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 442264 3340 442316 3392
rect 446220 3340 446272 3392
rect 449164 3340 449216 3392
rect 248788 3272 248840 3324
rect 324964 3272 325016 3324
rect 326804 3272 326856 3324
rect 31300 3204 31352 3256
rect 33784 3204 33836 3256
rect 143540 3204 143592 3256
rect 144828 3204 144880 3256
rect 168380 3204 168432 3256
rect 169668 3204 169720 3256
rect 173164 3204 173216 3256
rect 174544 3204 174596 3256
rect 222752 3204 222804 3256
rect 229744 3204 229796 3256
rect 242164 3204 242216 3256
rect 245200 3204 245252 3256
rect 250444 3204 250496 3256
rect 254676 3204 254728 3256
rect 385684 3204 385736 3256
rect 387156 3204 387208 3256
rect 485044 3340 485096 3392
rect 547880 3408 547932 3460
rect 558184 3408 558236 3460
rect 565636 3408 565688 3460
rect 490564 3340 490616 3392
rect 492312 3340 492364 3392
rect 497464 3340 497516 3392
rect 499396 3340 499448 3392
rect 515404 3340 515456 3392
rect 517152 3340 517204 3392
rect 465724 3272 465776 3324
rect 467472 3272 467524 3324
rect 482284 3272 482336 3324
rect 486424 3272 486476 3324
rect 500316 3272 500368 3324
rect 502984 3272 503036 3324
rect 580264 3272 580316 3324
rect 581000 3272 581052 3324
rect 458088 3204 458140 3256
rect 48964 3136 49016 3188
rect 53104 3136 53156 3188
rect 235816 3136 235868 3188
rect 238024 3136 238076 3188
rect 239312 3136 239364 3188
rect 240784 3136 240836 3188
rect 15936 3068 15988 3120
rect 201960 3068 202012 3120
rect 242532 3068 242584 3120
rect 247592 3068 247644 3120
rect 413284 3068 413336 3120
rect 420184 3068 420236 3120
rect 543004 3068 543056 3120
rect 545488 3068 545540 3120
rect 554044 3068 554096 3120
rect 556160 3068 556212 3120
rect 8760 3000 8812 3052
rect 14464 3000 14516 3052
rect 104532 3000 104584 3052
rect 105544 3000 105596 3052
rect 184940 3000 184992 3052
rect 187056 3000 187108 3052
rect 233424 3000 233476 3052
rect 234528 3000 234580 3052
rect 364984 3000 365036 3052
rect 367008 3000 367060 3052
rect 369124 3000 369176 3052
rect 371700 3000 371752 3052
rect 377404 3000 377456 3052
rect 379980 3000 380032 3052
rect 435364 3000 435416 3052
rect 437940 3000 437992 3052
rect 504364 3000 504416 3052
rect 510068 3000 510120 3052
rect 511264 3000 511316 3052
rect 513564 3000 513616 3052
rect 529204 3000 529256 3052
rect 531320 3000 531372 3052
rect 312544 2932 312596 2984
rect 315028 2932 315080 2984
rect 446404 2932 446456 2984
rect 452108 2932 452160 2984
rect 493324 2932 493376 2984
rect 495900 2932 495952 2984
rect 522304 2932 522356 2984
rect 524236 2932 524288 2984
rect 530676 2932 530728 2984
rect 532516 2932 532568 2984
rect 275284 2864 275336 2916
rect 279516 2864 279568 2916
rect 472716 2864 472768 2916
rect 474556 2864 474608 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 8128 700398 8156 703520
rect 24320 700466 24348 703520
rect 40512 700534 40540 703520
rect 72988 700602 73016 703520
rect 89180 700670 89208 703520
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 41328 700528 41380 700534
rect 41328 700470 41380 700476
rect 24308 700460 24360 700466
rect 24308 700402 24360 700408
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 670818 3464 671191
rect 3424 670812 3476 670818
rect 3424 670754 3476 670760
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 41340 327758 41368 700470
rect 105464 699718 105492 703520
rect 137848 700806 137876 703520
rect 154132 700874 154160 703520
rect 154120 700868 154172 700874
rect 154120 700810 154172 700816
rect 137836 700800 137888 700806
rect 137836 700742 137888 700748
rect 170324 699718 170352 703520
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 218992 700262 219020 703520
rect 218980 700256 219032 700262
rect 218980 700198 219032 700204
rect 235184 699718 235212 703520
rect 251180 701004 251232 701010
rect 251180 700946 251232 700952
rect 248328 700936 248380 700942
rect 248328 700878 248380 700884
rect 245568 700732 245620 700738
rect 245568 700674 245620 700680
rect 242808 700528 242860 700534
rect 242808 700470 242860 700476
rect 241336 700324 241388 700330
rect 241336 700266 241388 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 233148 699712 233200 699718
rect 233148 699654 233200 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 41328 327752 41380 327758
rect 41328 327694 41380 327700
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 106200 305862 106228 699654
rect 171060 305998 171088 699654
rect 231676 590708 231728 590714
rect 231676 590650 231728 590656
rect 198648 554192 198700 554198
rect 198648 554134 198700 554140
rect 198556 554056 198608 554062
rect 198556 553998 198608 554004
rect 198464 482316 198516 482322
rect 198464 482258 198516 482264
rect 171048 305992 171100 305998
rect 171048 305934 171100 305940
rect 106188 305856 106240 305862
rect 106188 305798 106240 305804
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 43444 303000 43496 303006
rect 43444 302942 43496 302948
rect 28264 302932 28316 302938
rect 28264 302874 28316 302880
rect 26884 302728 26936 302734
rect 26884 302670 26936 302676
rect 4804 302660 4856 302666
rect 4804 302602 4856 302608
rect 3884 298512 3936 298518
rect 3884 298454 3936 298460
rect 3424 298444 3476 298450
rect 3424 298386 3476 298392
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3436 241097 3464 298386
rect 3516 298376 3568 298382
rect 3516 298318 3568 298324
rect 3528 254153 3556 298318
rect 3896 293185 3924 298454
rect 3882 293176 3938 293185
rect 3882 293111 3938 293120
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4816 97782 4844 302602
rect 10324 301096 10376 301102
rect 10324 301038 10376 301044
rect 10336 267714 10364 301038
rect 11704 299804 11756 299810
rect 11704 299746 11756 299752
rect 10324 267708 10376 267714
rect 10324 267650 10376 267656
rect 11716 164218 11744 299746
rect 11704 164212 11756 164218
rect 11704 164154 11756 164160
rect 19248 98660 19300 98666
rect 19248 98602 19300 98608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 17868 95940 17920 95946
rect 17868 95882 17920 95888
rect 12346 94480 12402 94489
rect 12346 94415 12402 94424
rect 5448 86284 5500 86290
rect 5448 86226 5500 86232
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 5460 6914 5488 86226
rect 5276 6886 5488 6914
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 5276 480 5304 6886
rect 11152 3868 11204 3874
rect 11152 3810 11204 3816
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 3538
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8772 480 8800 2994
rect 9968 480 9996 3606
rect 11164 480 11192 3810
rect 12360 480 12388 94415
rect 14464 93152 14516 93158
rect 14464 93094 14516 93100
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13556 480 13584 3674
rect 14476 3058 14504 93094
rect 15844 87644 15896 87650
rect 15844 87586 15896 87592
rect 15856 3534 15884 87586
rect 17880 3602 17908 95882
rect 19260 3602 19288 98602
rect 25504 94512 25556 94518
rect 25504 94454 25556 94460
rect 23388 91792 23440 91798
rect 23388 91734 23440 91740
rect 21364 89004 21416 89010
rect 21364 88946 21416 88952
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14752 480 14780 3470
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 15948 480 15976 3062
rect 17052 480 17080 3538
rect 18248 480 18276 3538
rect 19444 480 19472 3946
rect 20628 3800 20680 3806
rect 20628 3742 20680 3748
rect 20640 480 20668 3742
rect 21376 3670 21404 88946
rect 23400 6914 23428 91734
rect 23032 6886 23428 6914
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21836 480 21864 3538
rect 23032 480 23060 6886
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24228 480 24256 5170
rect 25320 3664 25372 3670
rect 25320 3606 25372 3612
rect 25332 480 25360 3606
rect 25516 3602 25544 94454
rect 26516 7608 26568 7614
rect 26516 7550 26568 7556
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 26528 480 26556 7550
rect 26896 6866 26924 302670
rect 28276 202842 28304 302874
rect 29644 302864 29696 302870
rect 29644 302806 29696 302812
rect 28264 202836 28316 202842
rect 28264 202778 28316 202784
rect 29656 150414 29684 302806
rect 32404 302796 32456 302802
rect 32404 302738 32456 302744
rect 29644 150408 29696 150414
rect 29644 150350 29696 150356
rect 29644 98728 29696 98734
rect 29644 98670 29696 98676
rect 28264 86352 28316 86358
rect 28264 86294 28316 86300
rect 26884 6860 26936 6866
rect 26884 6802 26936 6808
rect 28276 3874 28304 86294
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 28264 3868 28316 3874
rect 28264 3810 28316 3816
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27724 480 27752 3538
rect 28920 480 28948 3878
rect 29656 3602 29684 98670
rect 32416 59362 32444 302738
rect 36544 98796 36596 98802
rect 36544 98738 36596 98744
rect 33784 94580 33836 94586
rect 33784 94522 33836 94528
rect 33048 86420 33100 86426
rect 33048 86362 33100 86368
rect 32404 59356 32456 59362
rect 32404 59298 32456 59304
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 29644 3596 29696 3602
rect 29644 3538 29696 3544
rect 30116 480 30144 8910
rect 33060 3602 33088 86362
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 31300 3256 31352 3262
rect 31300 3198 31352 3204
rect 31312 480 31340 3198
rect 32416 480 32444 3538
rect 33612 480 33640 8978
rect 33796 3262 33824 94522
rect 35164 89072 35216 89078
rect 35164 89014 35216 89020
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 33784 3256 33836 3262
rect 33784 3198 33836 3204
rect 34808 480 34836 4014
rect 35176 4010 35204 89014
rect 35992 5160 36044 5166
rect 35992 5102 36044 5108
rect 35164 4004 35216 4010
rect 35164 3946 35216 3952
rect 36004 480 36032 5102
rect 36556 3738 36584 98738
rect 39948 97300 40000 97306
rect 39948 97242 40000 97248
rect 39302 97200 39358 97209
rect 39302 97135 39358 97144
rect 37096 94648 37148 94654
rect 37096 94590 37148 94596
rect 37108 16574 37136 94590
rect 37108 16546 37228 16574
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 37200 480 37228 16546
rect 38384 6248 38436 6254
rect 38384 6190 38436 6196
rect 38396 480 38424 6190
rect 39316 3806 39344 97135
rect 39960 6914 39988 97242
rect 41328 90364 41380 90370
rect 41328 90306 41380 90312
rect 39592 6886 39988 6914
rect 39304 3800 39356 3806
rect 39304 3742 39356 3748
rect 39592 480 39620 6886
rect 41340 3602 41368 90306
rect 43456 20670 43484 302942
rect 152464 301300 152516 301306
rect 152464 301242 152516 301248
rect 148324 301164 148376 301170
rect 148324 301106 148376 301112
rect 101404 99272 101456 99278
rect 101404 99214 101456 99220
rect 94504 99204 94556 99210
rect 94504 99146 94556 99152
rect 93124 99136 93176 99142
rect 93124 99078 93176 99084
rect 71044 99068 71096 99074
rect 71044 99010 71096 99016
rect 57244 99000 57296 99006
rect 57244 98942 57296 98948
rect 50344 98932 50396 98938
rect 50344 98874 50396 98880
rect 46204 98864 46256 98870
rect 46204 98806 46256 98812
rect 45468 91860 45520 91866
rect 45468 91802 45520 91808
rect 44088 87712 44140 87718
rect 44088 87654 44140 87660
rect 43444 20664 43496 20670
rect 43444 20606 43496 20612
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 40696 480 40724 3538
rect 41892 480 41920 3674
rect 44100 3602 44128 87654
rect 45376 3800 45428 3806
rect 45376 3742 45428 3748
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 43088 480 43116 3538
rect 44284 480 44312 3538
rect 45388 1986 45416 3742
rect 45480 3602 45508 91802
rect 46216 4078 46244 98806
rect 47584 89140 47636 89146
rect 47584 89082 47636 89088
rect 46204 4072 46256 4078
rect 46204 4014 46256 4020
rect 47596 3942 47624 89082
rect 50160 7676 50212 7682
rect 50160 7618 50212 7624
rect 47860 5024 47912 5030
rect 47860 4966 47912 4972
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 46664 3868 46716 3874
rect 46664 3810 46716 3816
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45388 1958 45508 1986
rect 45480 480 45508 1958
rect 46676 480 46704 3810
rect 47872 480 47900 4966
rect 48964 3188 49016 3194
rect 48964 3130 49016 3136
rect 48976 480 49004 3130
rect 50172 480 50200 7618
rect 50356 3738 50384 98874
rect 54484 91928 54536 91934
rect 54484 91870 54536 91876
rect 53104 90432 53156 90438
rect 53104 90374 53156 90380
rect 50344 3732 50396 3738
rect 50344 3674 50396 3680
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 51368 480 51396 3674
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52564 480 52592 3538
rect 53116 3194 53144 90374
rect 53748 3936 53800 3942
rect 53748 3878 53800 3884
rect 53104 3188 53156 3194
rect 53104 3130 53156 3136
rect 53760 480 53788 3878
rect 54496 3602 54524 91870
rect 57256 6914 57284 98942
rect 58624 97368 58676 97374
rect 58624 97310 58676 97316
rect 57164 6886 57284 6914
rect 54944 5092 54996 5098
rect 54944 5034 54996 5040
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 54956 480 54984 5034
rect 56048 4004 56100 4010
rect 56048 3946 56100 3952
rect 56060 480 56088 3946
rect 57164 3806 57192 6886
rect 58636 5166 58664 97310
rect 70308 96008 70360 96014
rect 70308 95950 70360 95956
rect 64788 94716 64840 94722
rect 64788 94658 64840 94664
rect 62028 6316 62080 6322
rect 62028 6258 62080 6264
rect 58624 5160 58676 5166
rect 58624 5102 58676 5108
rect 58716 5160 58768 5166
rect 58716 5102 58768 5108
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57152 3800 57204 3806
rect 57152 3742 57204 3748
rect 57256 480 57284 4014
rect 58728 2666 58756 5102
rect 60832 4140 60884 4146
rect 60832 4082 60884 4088
rect 59636 3324 59688 3330
rect 59636 3266 59688 3272
rect 58452 2638 58756 2666
rect 58452 480 58480 2638
rect 59648 480 59676 3266
rect 60844 480 60872 4082
rect 62040 480 62068 6258
rect 63224 3800 63276 3806
rect 63224 3742 63276 3748
rect 63236 480 63264 3742
rect 64800 3602 64828 94658
rect 68284 93220 68336 93226
rect 68284 93162 68336 93168
rect 65524 90500 65576 90506
rect 65524 90442 65576 90448
rect 65536 4010 65564 90442
rect 65616 6384 65668 6390
rect 65616 6326 65668 6332
rect 65524 4004 65576 4010
rect 65524 3946 65576 3952
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 64340 480 64368 3538
rect 65628 3210 65656 6326
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 65536 3182 65656 3210
rect 65536 480 65564 3182
rect 66732 480 66760 3334
rect 67928 480 67956 3538
rect 68296 3330 68324 93162
rect 70216 89208 70268 89214
rect 70216 89150 70268 89156
rect 68928 47592 68980 47598
rect 68928 47534 68980 47540
rect 68940 3602 68968 47534
rect 70228 16574 70256 89150
rect 70136 16546 70256 16574
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 68284 3324 68336 3330
rect 68284 3266 68336 3272
rect 69124 480 69152 3538
rect 70136 3482 70164 16546
rect 70320 6914 70348 95950
rect 70228 6886 70348 6914
rect 70228 3602 70256 6886
rect 71056 4146 71084 99010
rect 78588 94784 78640 94790
rect 78588 94726 78640 94732
rect 73068 93288 73120 93294
rect 73068 93230 73120 93236
rect 71044 4140 71096 4146
rect 71044 4082 71096 4088
rect 71504 4004 71556 4010
rect 71504 3946 71556 3952
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 70136 3454 70348 3482
rect 70320 480 70348 3454
rect 71516 480 71544 3946
rect 73080 3602 73108 93230
rect 77208 91996 77260 92002
rect 77208 91938 77260 91944
rect 75184 90568 75236 90574
rect 75184 90510 75236 90516
rect 75000 7948 75052 7954
rect 75000 7890 75052 7896
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 72608 3596 72660 3602
rect 72608 3538 72660 3544
rect 73068 3596 73120 3602
rect 73068 3538 73120 3544
rect 72620 480 72648 3538
rect 73816 480 73844 4082
rect 75012 480 75040 7890
rect 75196 3398 75224 90510
rect 77220 3602 77248 91938
rect 76196 3596 76248 3602
rect 76196 3538 76248 3544
rect 77208 3596 77260 3602
rect 77208 3538 77260 3544
rect 77392 3596 77444 3602
rect 77392 3538 77444 3544
rect 75184 3392 75236 3398
rect 75184 3334 75236 3340
rect 76208 480 76236 3538
rect 77404 480 77432 3538
rect 78600 480 78628 94726
rect 84108 93356 84160 93362
rect 84108 93298 84160 93304
rect 79968 92064 80020 92070
rect 79968 92006 80020 92012
rect 79324 89276 79376 89282
rect 79324 89218 79376 89224
rect 79336 3602 79364 89218
rect 79980 6914 80008 92006
rect 80704 89344 80756 89350
rect 80704 89286 80756 89292
rect 79704 6886 80008 6914
rect 79324 3596 79376 3602
rect 79324 3538 79376 3544
rect 79704 480 79732 6886
rect 80716 4146 80744 89286
rect 80704 4140 80756 4146
rect 80704 4082 80756 4088
rect 82084 4140 82136 4146
rect 82084 4082 82136 4088
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 80900 480 80928 3334
rect 82096 480 82124 4082
rect 84120 3602 84148 93298
rect 90364 90636 90416 90642
rect 90364 90578 90416 90584
rect 88984 87916 89036 87922
rect 88984 87858 89036 87864
rect 87604 87848 87656 87854
rect 87604 87790 87656 87796
rect 86224 87780 86276 87786
rect 86224 87722 86276 87728
rect 85488 10328 85540 10334
rect 85488 10270 85540 10276
rect 85500 3602 85528 10270
rect 85672 6452 85724 6458
rect 85672 6394 85724 6400
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 84108 3596 84160 3602
rect 84108 3538 84160 3544
rect 84476 3596 84528 3602
rect 84476 3538 84528 3544
rect 85488 3596 85540 3602
rect 85488 3538 85540 3544
rect 83292 480 83320 3538
rect 84488 480 84516 3538
rect 85684 480 85712 6394
rect 86236 3398 86264 87722
rect 86868 9104 86920 9110
rect 86868 9046 86920 9052
rect 86224 3392 86276 3398
rect 86224 3334 86276 3340
rect 86880 480 86908 9046
rect 87616 4078 87644 87790
rect 87972 10396 88024 10402
rect 87972 10338 88024 10344
rect 87604 4072 87656 4078
rect 87604 4014 87656 4020
rect 87984 480 88012 10338
rect 88996 3942 89024 87858
rect 88984 3936 89036 3942
rect 88984 3878 89036 3884
rect 90376 3602 90404 90578
rect 92388 10464 92440 10470
rect 92388 10406 92440 10412
rect 90456 9172 90508 9178
rect 90456 9114 90508 9120
rect 89168 3596 89220 3602
rect 89168 3538 89220 3544
rect 90364 3596 90416 3602
rect 90364 3538 90416 3544
rect 89180 480 89208 3538
rect 90468 3482 90496 9114
rect 92400 3602 92428 10406
rect 93136 4146 93164 99078
rect 93952 9240 94004 9246
rect 93952 9182 94004 9188
rect 93124 4140 93176 4146
rect 93124 4082 93176 4088
rect 92756 3936 92808 3942
rect 92756 3878 92808 3884
rect 91560 3596 91612 3602
rect 91560 3538 91612 3544
rect 92388 3596 92440 3602
rect 92388 3538 92440 3544
rect 90376 3454 90496 3482
rect 90376 480 90404 3454
rect 91572 480 91600 3538
rect 92768 480 92796 3878
rect 93964 480 93992 9182
rect 94516 3874 94544 99146
rect 97264 97436 97316 97442
rect 97264 97378 97316 97384
rect 95148 10532 95200 10538
rect 95148 10474 95200 10480
rect 94504 3868 94556 3874
rect 94504 3810 94556 3816
rect 95160 480 95188 10474
rect 97276 3942 97304 97378
rect 98644 96824 98696 96830
rect 98644 96766 98696 96772
rect 97448 9308 97500 9314
rect 97448 9250 97500 9256
rect 97264 3936 97316 3942
rect 97264 3878 97316 3884
rect 96252 3868 96304 3874
rect 96252 3810 96304 3816
rect 96264 480 96292 3810
rect 97460 480 97488 9250
rect 98656 5234 98684 96766
rect 99288 10600 99340 10606
rect 99288 10542 99340 10548
rect 98644 5228 98696 5234
rect 98644 5170 98696 5176
rect 99300 3602 99328 10542
rect 99840 5228 99892 5234
rect 99840 5170 99892 5176
rect 98644 3596 98696 3602
rect 98644 3538 98696 3544
rect 99288 3596 99340 3602
rect 99288 3538 99340 3544
rect 98656 480 98684 3538
rect 99852 480 99880 5170
rect 101036 4072 101088 4078
rect 101036 4014 101088 4020
rect 101048 480 101076 4014
rect 101416 4010 101444 99214
rect 134524 97912 134576 97918
rect 134524 97854 134576 97860
rect 126888 97844 126940 97850
rect 126888 97786 126940 97792
rect 124864 97776 124916 97782
rect 124864 97718 124916 97724
rect 119344 97640 119396 97646
rect 119344 97582 119396 97588
rect 115204 97572 115256 97578
rect 115204 97514 115256 97520
rect 104164 92132 104216 92138
rect 104164 92074 104216 92080
rect 103428 89412 103480 89418
rect 103428 89354 103480 89360
rect 101404 4004 101456 4010
rect 101404 3946 101456 3952
rect 103336 4004 103388 4010
rect 103336 3946 103388 3952
rect 102232 3596 102284 3602
rect 102232 3538 102284 3544
rect 102244 480 102272 3538
rect 103348 480 103376 3946
rect 103440 3602 103468 89354
rect 104176 4078 104204 92074
rect 112444 90840 112496 90846
rect 112444 90782 112496 90788
rect 108948 90772 109000 90778
rect 108948 90714 109000 90720
rect 105544 90704 105596 90710
rect 105544 90646 105596 90652
rect 104164 4072 104216 4078
rect 104164 4014 104216 4020
rect 103428 3596 103480 3602
rect 103428 3538 103480 3544
rect 105556 3058 105584 90646
rect 107568 84856 107620 84862
rect 107568 84798 107620 84804
rect 106188 15904 106240 15910
rect 106188 15846 106240 15852
rect 106200 3602 106228 15846
rect 107580 3602 107608 84798
rect 108960 3602 108988 90714
rect 111064 87984 111116 87990
rect 111064 87926 111116 87932
rect 111076 3602 111104 87926
rect 111708 11756 111760 11762
rect 111708 11698 111760 11704
rect 105728 3596 105780 3602
rect 105728 3538 105780 3544
rect 106188 3596 106240 3602
rect 106188 3538 106240 3544
rect 106924 3596 106976 3602
rect 106924 3538 106976 3544
rect 107568 3596 107620 3602
rect 107568 3538 107620 3544
rect 108120 3596 108172 3602
rect 108120 3538 108172 3544
rect 108948 3596 109000 3602
rect 108948 3538 109000 3544
rect 109316 3596 109368 3602
rect 109316 3538 109368 3544
rect 111064 3596 111116 3602
rect 111064 3538 111116 3544
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 104532 3052 104584 3058
rect 104532 2994 104584 3000
rect 105544 3052 105596 3058
rect 105544 2994 105596 3000
rect 104544 480 104572 2994
rect 105740 480 105768 3538
rect 106936 480 106964 3538
rect 108132 480 108160 3538
rect 109328 480 109356 3538
rect 110512 3392 110564 3398
rect 110512 3334 110564 3340
rect 110524 480 110552 3334
rect 111628 480 111656 3538
rect 111720 3398 111748 11698
rect 112456 3602 112484 90782
rect 112812 3936 112864 3942
rect 112812 3878 112864 3884
rect 112444 3596 112496 3602
rect 112444 3538 112496 3544
rect 111708 3392 111760 3398
rect 111708 3334 111760 3340
rect 112824 480 112852 3878
rect 115216 3602 115244 97514
rect 116584 89480 116636 89486
rect 116584 89422 116636 89428
rect 115296 9376 115348 9382
rect 115296 9318 115348 9324
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 114020 480 114048 3538
rect 115308 3482 115336 9318
rect 116596 3942 116624 89422
rect 119356 11762 119384 97582
rect 124128 89548 124180 89554
rect 124128 89490 124180 89496
rect 122104 86488 122156 86494
rect 122104 86430 122156 86436
rect 119344 11756 119396 11762
rect 119344 11698 119396 11704
rect 119896 11756 119948 11762
rect 119896 11698 119948 11704
rect 117228 10668 117280 10674
rect 117228 10610 117280 10616
rect 116584 3936 116636 3942
rect 116584 3878 116636 3884
rect 117240 3602 117268 10610
rect 118792 9444 118844 9450
rect 118792 9386 118844 9392
rect 117596 4004 117648 4010
rect 117596 3946 117648 3952
rect 116400 3596 116452 3602
rect 116400 3538 116452 3544
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 115216 3454 115336 3482
rect 115216 480 115244 3454
rect 116412 480 116440 3538
rect 117608 480 117636 3946
rect 118804 480 118832 9386
rect 119908 480 119936 11698
rect 122116 4078 122144 86430
rect 122288 9512 122340 9518
rect 122288 9454 122340 9460
rect 122104 4072 122156 4078
rect 122104 4014 122156 4020
rect 121092 3936 121144 3942
rect 121092 3878 121144 3884
rect 121104 480 121132 3878
rect 122300 480 122328 9454
rect 124140 3602 124168 89490
rect 124876 5302 124904 97718
rect 126244 97708 126296 97714
rect 126244 97650 126296 97656
rect 124864 5296 124916 5302
rect 124864 5238 124916 5244
rect 126256 4214 126284 97650
rect 124680 4208 124732 4214
rect 124680 4150 124732 4156
rect 126244 4208 126296 4214
rect 126244 4150 126296 4156
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 123496 480 123524 3538
rect 124692 480 124720 4150
rect 126900 3602 126928 97786
rect 133788 96076 133840 96082
rect 133788 96018 133840 96024
rect 128268 94852 128320 94858
rect 128268 94794 128320 94800
rect 128176 92200 128228 92206
rect 128176 92142 128228 92148
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 126888 3596 126940 3602
rect 126888 3538 126940 3544
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 125888 480 125916 3538
rect 126992 480 127020 3538
rect 128188 480 128216 92142
rect 128280 3602 128308 94794
rect 131028 93424 131080 93430
rect 131028 93366 131080 93372
rect 129372 4072 129424 4078
rect 129372 4014 129424 4020
rect 128268 3596 128320 3602
rect 128268 3538 128320 3544
rect 129384 480 129412 4014
rect 131040 3602 131068 93366
rect 131764 7744 131816 7750
rect 131764 7686 131816 7692
rect 130568 3596 130620 3602
rect 130568 3538 130620 3544
rect 131028 3596 131080 3602
rect 131028 3538 131080 3544
rect 130580 480 130608 3538
rect 131776 480 131804 7686
rect 133800 3602 133828 96018
rect 134156 6520 134208 6526
rect 134156 6462 134208 6468
rect 132960 3596 133012 3602
rect 132960 3538 133012 3544
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 132972 480 133000 3538
rect 134168 480 134196 6462
rect 134536 6458 134564 97854
rect 142804 97232 142856 97238
rect 142804 97174 142856 97180
rect 137284 94920 137336 94926
rect 137284 94862 137336 94868
rect 135260 7540 135312 7546
rect 135260 7482 135312 7488
rect 134524 6452 134576 6458
rect 134524 6394 134576 6400
rect 135272 480 135300 7482
rect 137296 3602 137324 94862
rect 142068 93492 142120 93498
rect 142068 93434 142120 93440
rect 138848 7812 138900 7818
rect 138848 7754 138900 7760
rect 137652 6520 137704 6526
rect 137652 6462 137704 6468
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 137284 3596 137336 3602
rect 137284 3538 137336 3544
rect 136468 480 136496 3538
rect 137664 480 137692 6462
rect 138860 480 138888 7754
rect 140044 3596 140096 3602
rect 140044 3538 140096 3544
rect 140056 480 140084 3538
rect 142080 3398 142108 93434
rect 142816 8022 142844 97174
rect 144828 95056 144880 95062
rect 144828 94998 144880 95004
rect 144736 93560 144788 93566
rect 144736 93502 144788 93508
rect 142804 8016 142856 8022
rect 142804 7958 142856 7964
rect 142436 7948 142488 7954
rect 142436 7890 142488 7896
rect 141240 3392 141292 3398
rect 141240 3334 141292 3340
rect 142068 3392 142120 3398
rect 142068 3334 142120 3340
rect 141252 480 141280 3334
rect 142448 480 142476 7890
rect 143540 3256 143592 3262
rect 143540 3198 143592 3204
rect 143552 480 143580 3198
rect 144748 480 144776 93502
rect 144840 3262 144868 94998
rect 147588 94988 147640 94994
rect 147588 94930 147640 94936
rect 146208 90908 146260 90914
rect 146208 90850 146260 90856
rect 146220 6914 146248 90850
rect 146944 7812 146996 7818
rect 146944 7754 146996 7760
rect 146956 7546 146984 7754
rect 146944 7540 146996 7546
rect 146944 7482 146996 7488
rect 145944 6886 146248 6914
rect 144828 3256 144880 3262
rect 144828 3198 144880 3204
rect 145944 480 145972 6886
rect 146944 4140 146996 4146
rect 146944 4082 146996 4088
rect 146956 3602 146984 4082
rect 147600 3602 147628 94930
rect 148336 45558 148364 301106
rect 151084 299872 151136 299878
rect 151084 299814 151136 299820
rect 150348 97980 150400 97986
rect 150348 97922 150400 97928
rect 148968 93696 149020 93702
rect 148968 93638 149020 93644
rect 148324 45552 148376 45558
rect 148324 45494 148376 45500
rect 148980 3602 149008 93638
rect 150360 3602 150388 97922
rect 151096 85542 151124 299814
rect 152476 137970 152504 301242
rect 156604 301232 156656 301238
rect 156604 301174 156656 301180
rect 155224 300076 155276 300082
rect 155224 300018 155276 300024
rect 155236 189038 155264 300018
rect 155224 189032 155276 189038
rect 155224 188974 155276 188980
rect 152464 137964 152516 137970
rect 152464 137906 152516 137912
rect 155224 96144 155276 96150
rect 155224 96086 155276 96092
rect 153108 93628 153160 93634
rect 153108 93570 153160 93576
rect 153016 90976 153068 90982
rect 153016 90918 153068 90924
rect 151084 85536 151136 85542
rect 151084 85478 151136 85484
rect 146944 3596 146996 3602
rect 146944 3538 146996 3544
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 147588 3596 147640 3602
rect 147588 3538 147640 3544
rect 148324 3596 148376 3602
rect 148324 3538 148376 3544
rect 148968 3596 149020 3602
rect 148968 3538 149020 3544
rect 149520 3596 149572 3602
rect 149520 3538 149572 3544
rect 150348 3596 150400 3602
rect 150348 3538 150400 3544
rect 151820 3596 151872 3602
rect 151820 3538 151872 3544
rect 147140 480 147168 3538
rect 148336 480 148364 3538
rect 149532 480 149560 3538
rect 150624 3392 150676 3398
rect 150624 3334 150676 3340
rect 150636 480 150664 3334
rect 151832 480 151860 3538
rect 153028 480 153056 90918
rect 153120 3602 153148 93570
rect 155236 3602 155264 96086
rect 155868 93764 155920 93770
rect 155868 93706 155920 93712
rect 155880 3602 155908 93706
rect 156616 33114 156644 301174
rect 159364 300008 159416 300014
rect 159364 299950 159416 299956
rect 157984 299940 158036 299946
rect 157984 299882 158036 299888
rect 157248 94376 157300 94382
rect 157248 94318 157300 94324
rect 156604 33108 156656 33114
rect 156604 33050 156656 33056
rect 157260 3602 157288 94318
rect 157996 71738 158024 299882
rect 159376 111790 159404 299950
rect 198476 298897 198504 482258
rect 198462 298888 198518 298897
rect 198462 298823 198518 298832
rect 198464 298580 198516 298586
rect 198464 298522 198516 298528
rect 198476 294681 198504 298522
rect 198568 296857 198596 553998
rect 198554 296848 198610 296857
rect 198554 296783 198610 296792
rect 198462 294672 198518 294681
rect 198462 294607 198518 294616
rect 198660 292641 198688 554134
rect 230388 536852 230440 536858
rect 230388 536794 230440 536800
rect 230296 524476 230348 524482
rect 230296 524418 230348 524424
rect 227628 470620 227680 470626
rect 227628 470562 227680 470568
rect 226156 456816 226208 456822
rect 226156 456758 226208 456764
rect 223396 404388 223448 404394
rect 223396 404330 223448 404336
rect 222108 378208 222160 378214
rect 222108 378150 222160 378156
rect 219348 324352 219400 324358
rect 219348 324294 219400 324300
rect 212172 303204 212224 303210
rect 212172 303146 212224 303152
rect 207112 303136 207164 303142
rect 207112 303078 207164 303084
rect 204628 303068 204680 303074
rect 204628 303010 204680 303016
rect 202052 302456 202104 302462
rect 202052 302398 202104 302404
rect 199384 301640 199436 301646
rect 199384 301582 199436 301588
rect 198646 292632 198702 292641
rect 198646 292567 198702 292576
rect 197358 290456 197414 290465
rect 197358 290391 197414 290400
rect 197372 289882 197400 290391
rect 170404 289876 170456 289882
rect 170404 289818 170456 289824
rect 197360 289876 197412 289882
rect 197360 289818 197412 289824
rect 160100 281580 160152 281586
rect 160100 281522 160152 281528
rect 160112 171134 160140 281522
rect 160112 171106 160600 171134
rect 160572 160698 160600 171106
rect 169208 160744 169260 160750
rect 160572 160670 160954 160698
rect 168958 160692 169208 160698
rect 168958 160686 169260 160692
rect 168958 160670 169248 160686
rect 162872 158574 162900 160004
rect 164896 158642 164924 160004
rect 166920 158710 166948 160004
rect 170416 158710 170444 289818
rect 198554 288416 198610 288425
rect 198554 288351 198610 288360
rect 198568 287094 198596 288351
rect 178684 287088 178736 287094
rect 178684 287030 178736 287036
rect 198556 287088 198608 287094
rect 198556 287030 198608 287036
rect 174544 282940 174596 282946
rect 174544 282882 174596 282888
rect 171784 242956 171836 242962
rect 171784 242898 171836 242904
rect 170496 222896 170548 222902
rect 170496 222838 170548 222844
rect 166908 158704 166960 158710
rect 166908 158646 166960 158652
rect 170404 158704 170456 158710
rect 170404 158646 170456 158652
rect 170508 158642 170536 222838
rect 171140 179240 171192 179246
rect 171138 179208 171140 179217
rect 171192 179208 171194 179217
rect 171138 179143 171194 179152
rect 171796 170513 171824 242898
rect 171876 238808 171928 238814
rect 171876 238750 171928 238756
rect 171782 170504 171838 170513
rect 171782 170439 171838 170448
rect 171888 168201 171916 238750
rect 171968 234660 172020 234666
rect 171968 234602 172020 234608
rect 171874 168192 171930 168201
rect 171874 168127 171930 168136
rect 171980 164529 172008 234602
rect 172060 233300 172112 233306
rect 172060 233242 172112 233248
rect 171966 164520 172022 164529
rect 171966 164455 172022 164464
rect 172072 164121 172100 233242
rect 173256 202904 173308 202910
rect 173256 202846 173308 202852
rect 173164 201544 173216 201550
rect 173164 201486 173216 201492
rect 172428 190120 172480 190126
rect 172428 190062 172480 190068
rect 172440 189961 172468 190062
rect 172426 189952 172482 189961
rect 172426 189887 172482 189896
rect 172428 189032 172480 189038
rect 172428 188974 172480 188980
rect 172440 188737 172468 188974
rect 172426 188728 172482 188737
rect 172426 188663 172482 188672
rect 172428 187672 172480 187678
rect 172428 187614 172480 187620
rect 172440 187377 172468 187614
rect 172426 187368 172482 187377
rect 172426 187303 172482 187312
rect 172428 186244 172480 186250
rect 172428 186186 172480 186192
rect 172440 186153 172468 186186
rect 172426 186144 172482 186153
rect 172426 186079 172482 186088
rect 172336 184884 172388 184890
rect 172336 184826 172388 184832
rect 172348 184385 172376 184826
rect 172428 184816 172480 184822
rect 172426 184784 172428 184793
rect 172480 184784 172482 184793
rect 172426 184719 172482 184728
rect 172334 184376 172390 184385
rect 172334 184311 172390 184320
rect 172428 183524 172480 183530
rect 172428 183466 172480 183472
rect 172440 183025 172468 183466
rect 172426 183016 172482 183025
rect 172426 182951 172482 182960
rect 172428 182164 172480 182170
rect 172428 182106 172480 182112
rect 172440 181801 172468 182106
rect 172426 181792 172482 181801
rect 172426 181727 172482 181736
rect 172428 180804 172480 180810
rect 172428 180746 172480 180752
rect 172440 180577 172468 180746
rect 172426 180568 172482 180577
rect 172426 180503 172482 180512
rect 172244 178016 172296 178022
rect 172244 177958 172296 177964
rect 172426 177984 172482 177993
rect 172256 177449 172284 177958
rect 172426 177919 172428 177928
rect 172480 177919 172482 177928
rect 172428 177890 172480 177896
rect 172242 177440 172298 177449
rect 172242 177375 172298 177384
rect 172244 176656 172296 176662
rect 172244 176598 172296 176604
rect 172256 176089 172284 176598
rect 172242 176080 172298 176089
rect 172242 176015 172298 176024
rect 172428 175228 172480 175234
rect 172428 175170 172480 175176
rect 172440 174865 172468 175170
rect 172426 174856 172482 174865
rect 172426 174791 172482 174800
rect 172428 173868 172480 173874
rect 172428 173810 172480 173816
rect 172440 173641 172468 173810
rect 172426 173632 172482 173641
rect 172426 173567 172482 173576
rect 172428 172440 172480 172446
rect 172426 172408 172428 172417
rect 172480 172408 172482 172417
rect 172426 172343 172482 172352
rect 172428 171080 172480 171086
rect 172426 171048 172428 171057
rect 172480 171048 172482 171057
rect 172426 170983 172482 170992
rect 172244 169720 172296 169726
rect 172244 169662 172296 169668
rect 172256 169153 172284 169662
rect 172242 169144 172298 169153
rect 172242 169079 172298 169088
rect 172428 167000 172480 167006
rect 172428 166942 172480 166948
rect 172440 166705 172468 166942
rect 172426 166696 172482 166705
rect 172426 166631 172482 166640
rect 172152 165572 172204 165578
rect 172152 165514 172204 165520
rect 172058 164112 172114 164121
rect 172058 164047 172114 164056
rect 171784 163668 171836 163674
rect 171784 163610 171836 163616
rect 164884 158636 164936 158642
rect 164884 158578 164936 158584
rect 170496 158636 170548 158642
rect 170496 158578 170548 158584
rect 162860 158568 162912 158574
rect 162860 158510 162912 158516
rect 171692 151768 171744 151774
rect 171692 151710 171744 151716
rect 171704 151609 171732 151710
rect 171690 151600 171746 151609
rect 171690 151535 171746 151544
rect 171508 151496 171560 151502
rect 171508 151438 171560 151444
rect 171520 151065 171548 151438
rect 171506 151056 171562 151065
rect 171506 150991 171562 151000
rect 171600 150612 171652 150618
rect 171600 150554 171652 150560
rect 171612 150521 171640 150554
rect 171598 150512 171654 150521
rect 171598 150447 171654 150456
rect 171692 150408 171744 150414
rect 171692 150350 171744 150356
rect 171704 149977 171732 150350
rect 171690 149968 171746 149977
rect 171690 149903 171746 149912
rect 171692 149456 171744 149462
rect 171690 149424 171692 149433
rect 171744 149424 171746 149433
rect 171690 149359 171746 149368
rect 171692 148844 171744 148850
rect 171692 148786 171744 148792
rect 171704 148345 171732 148786
rect 171690 148336 171746 148345
rect 171690 148271 171746 148280
rect 171508 147892 171560 147898
rect 171508 147834 171560 147840
rect 171520 147801 171548 147834
rect 171506 147792 171562 147801
rect 171506 147727 171562 147736
rect 171508 147552 171560 147558
rect 171508 147494 171560 147500
rect 171520 146713 171548 147494
rect 171506 146704 171562 146713
rect 171506 146639 171562 146648
rect 171508 145852 171560 145858
rect 171508 145794 171560 145800
rect 171520 145081 171548 145794
rect 171506 145072 171562 145081
rect 171506 145007 171562 145016
rect 171600 144220 171652 144226
rect 171600 144162 171652 144168
rect 171508 142860 171560 142866
rect 171508 142802 171560 142808
rect 171416 141976 171468 141982
rect 171414 141944 171416 141953
rect 171468 141944 171470 141953
rect 171414 141879 171470 141888
rect 171520 141409 171548 142802
rect 171612 142497 171640 144162
rect 171796 144129 171824 163610
rect 172164 162353 172192 165514
rect 172244 164212 172296 164218
rect 172244 164154 172296 164160
rect 172256 163577 172284 164154
rect 172242 163568 172298 163577
rect 172242 163503 172298 163512
rect 172150 162344 172206 162353
rect 172150 162279 172206 162288
rect 172428 161288 172480 161294
rect 172428 161230 172480 161236
rect 172440 160993 172468 161230
rect 172426 160984 172482 160993
rect 172426 160919 172482 160928
rect 171968 156664 172020 156670
rect 171968 156606 172020 156612
rect 171782 144120 171838 144129
rect 171782 144055 171838 144064
rect 171980 143585 172008 156606
rect 172336 154556 172388 154562
rect 172336 154498 172388 154504
rect 172244 154488 172296 154494
rect 172244 154430 172296 154436
rect 172256 153241 172284 154430
rect 172348 153785 172376 154498
rect 172334 153776 172390 153785
rect 172334 153711 172390 153720
rect 172242 153232 172298 153241
rect 172242 153167 172298 153176
rect 172428 153196 172480 153202
rect 172428 153138 172480 153144
rect 172336 153128 172388 153134
rect 172336 153070 172388 153076
rect 172348 152153 172376 153070
rect 172440 152697 172468 153138
rect 172426 152688 172482 152697
rect 172426 152623 172482 152632
rect 172334 152144 172390 152153
rect 172334 152079 172390 152088
rect 173176 150414 173204 201486
rect 173268 150618 173296 202846
rect 173440 198756 173492 198762
rect 173440 198698 173492 198704
rect 173348 197396 173400 197402
rect 173348 197338 173400 197344
rect 173256 150612 173308 150618
rect 173256 150554 173308 150560
rect 173164 150408 173216 150414
rect 173164 150350 173216 150356
rect 173360 148918 173388 197338
rect 173452 149462 173480 198698
rect 173532 194608 173584 194614
rect 173532 194550 173584 194556
rect 173440 149456 173492 149462
rect 173440 149398 173492 149404
rect 172244 148912 172296 148918
rect 172242 148880 172244 148889
rect 173348 148912 173400 148918
rect 172296 148880 172298 148889
rect 173348 148854 173400 148860
rect 173544 148850 173572 194550
rect 173624 193248 173676 193254
rect 173624 193190 173676 193196
rect 172242 148815 172298 148824
rect 173532 148844 173584 148850
rect 173532 148786 173584 148792
rect 173164 148368 173216 148374
rect 173164 148310 173216 148316
rect 172428 147620 172480 147626
rect 172428 147562 172480 147568
rect 172440 147257 172468 147562
rect 172426 147248 172482 147257
rect 172426 147183 172482 147192
rect 172428 146260 172480 146266
rect 172428 146202 172480 146208
rect 172336 146192 172388 146198
rect 172334 146160 172336 146169
rect 172388 146160 172390 146169
rect 172334 146095 172390 146104
rect 172440 145625 172468 146202
rect 172426 145616 172482 145625
rect 172426 145551 172482 145560
rect 172428 144900 172480 144906
rect 172428 144842 172480 144848
rect 172440 144537 172468 144842
rect 172426 144528 172482 144537
rect 172426 144463 172482 144472
rect 171966 143576 172022 143585
rect 171966 143511 172022 143520
rect 172244 143540 172296 143546
rect 172244 143482 172296 143488
rect 172256 143041 172284 143482
rect 172242 143032 172298 143041
rect 172242 142967 172298 142976
rect 171598 142488 171654 142497
rect 171598 142423 171654 142432
rect 172428 142112 172480 142118
rect 172428 142054 172480 142060
rect 171506 141400 171562 141409
rect 171506 141335 171562 141344
rect 171508 141296 171560 141302
rect 171508 141238 171560 141244
rect 171520 140321 171548 141238
rect 172440 140865 172468 142054
rect 172426 140856 172482 140865
rect 172426 140791 172482 140800
rect 171506 140312 171562 140321
rect 171506 140247 171562 140256
rect 172244 140072 172296 140078
rect 172244 140014 172296 140020
rect 171692 139800 171744 139806
rect 171690 139768 171692 139777
rect 171744 139768 171746 139777
rect 171690 139703 171746 139712
rect 171876 138916 171928 138922
rect 171876 138858 171928 138864
rect 171692 138780 171744 138786
rect 171692 138722 171744 138728
rect 171704 138145 171732 138722
rect 171888 138689 171916 138858
rect 171874 138680 171930 138689
rect 171874 138615 171930 138624
rect 171690 138136 171746 138145
rect 171690 138071 171746 138080
rect 172256 137057 172284 140014
rect 173176 139806 173204 148310
rect 173636 147898 173664 193190
rect 174556 158574 174584 282882
rect 175924 278792 175976 278798
rect 175924 278734 175976 278740
rect 174636 229152 174688 229158
rect 174636 229094 174688 229100
rect 174648 165578 174676 229094
rect 175936 190126 175964 278734
rect 177396 247104 177448 247110
rect 177396 247046 177448 247052
rect 176016 226364 176068 226370
rect 176016 226306 176068 226312
rect 175924 190120 175976 190126
rect 175924 190062 175976 190068
rect 174728 186380 174780 186386
rect 174728 186322 174780 186328
rect 174636 165572 174688 165578
rect 174636 165514 174688 165520
rect 174544 158568 174596 158574
rect 174544 158510 174596 158516
rect 174544 154624 174596 154630
rect 174544 154566 174596 154572
rect 173624 147892 173676 147898
rect 173624 147834 173676 147840
rect 173164 139800 173216 139806
rect 173164 139742 173216 139748
rect 172428 139324 172480 139330
rect 172428 139266 172480 139272
rect 172440 139233 172468 139266
rect 172426 139224 172482 139233
rect 172426 139159 172482 139168
rect 174556 138786 174584 154566
rect 174740 146198 174768 186322
rect 176028 161294 176056 226306
rect 177304 225004 177356 225010
rect 177304 224946 177356 224952
rect 176108 189100 176160 189106
rect 176108 189042 176160 189048
rect 176016 161288 176068 161294
rect 176016 161230 176068 161236
rect 175924 157412 175976 157418
rect 175924 157354 175976 157360
rect 174728 146192 174780 146198
rect 174728 146134 174780 146140
rect 175936 138922 175964 157354
rect 176120 147558 176148 189042
rect 176108 147552 176160 147558
rect 176108 147494 176160 147500
rect 175924 138916 175976 138922
rect 175924 138858 175976 138864
rect 174544 138780 174596 138786
rect 174544 138722 174596 138728
rect 175924 138032 175976 138038
rect 175924 137974 175976 137980
rect 172428 137964 172480 137970
rect 172428 137906 172480 137912
rect 172440 137601 172468 137906
rect 172426 137592 172482 137601
rect 172426 137527 172482 137536
rect 172336 137284 172388 137290
rect 172336 137226 172388 137232
rect 172242 137048 172298 137057
rect 172242 136983 172298 136992
rect 172244 136536 172296 136542
rect 172348 136513 172376 137226
rect 172520 136672 172572 136678
rect 172520 136614 172572 136620
rect 172428 136604 172480 136610
rect 172428 136546 172480 136552
rect 172244 136478 172296 136484
rect 172334 136504 172390 136513
rect 170404 135924 170456 135930
rect 170404 135866 170456 135872
rect 160940 122874 160968 124100
rect 160928 122868 160980 122874
rect 160928 122810 160980 122816
rect 162872 122738 162900 124100
rect 164896 122806 164924 124100
rect 164884 122800 164936 122806
rect 164884 122742 164936 122748
rect 162860 122732 162912 122738
rect 162860 122674 162912 122680
rect 159364 111784 159416 111790
rect 159364 111726 159416 111732
rect 166920 99414 166948 124100
rect 168944 122942 168972 124100
rect 168932 122936 168984 122942
rect 168932 122878 168984 122884
rect 170416 122806 170444 135866
rect 172256 135425 172284 136478
rect 172334 136439 172390 136448
rect 172440 135969 172468 136546
rect 172426 135960 172482 135969
rect 172426 135895 172482 135904
rect 172242 135416 172298 135425
rect 172242 135351 172298 135360
rect 172244 135312 172296 135318
rect 172244 135254 172296 135260
rect 171692 135244 171744 135250
rect 171692 135186 171744 135192
rect 171704 133929 171732 135186
rect 171876 135176 171928 135182
rect 171876 135118 171928 135124
rect 171888 134337 171916 135118
rect 172256 134881 172284 135254
rect 172242 134872 172298 134881
rect 172242 134807 172298 134816
rect 171874 134328 171930 134337
rect 171874 134263 171930 134272
rect 172428 133952 172480 133958
rect 171690 133920 171746 133929
rect 172428 133894 172480 133900
rect 171690 133855 171746 133864
rect 172440 132841 172468 133894
rect 172532 133385 172560 136614
rect 175936 135250 175964 137974
rect 175924 135244 175976 135250
rect 175924 135186 175976 135192
rect 172518 133376 172574 133385
rect 172518 133311 172574 133320
rect 172426 132832 172482 132841
rect 172426 132767 172482 132776
rect 171140 132524 171192 132530
rect 171140 132466 171192 132472
rect 171152 132297 171180 132466
rect 171138 132288 171194 132297
rect 171138 132223 171194 132232
rect 172426 131744 172482 131753
rect 172426 131679 172482 131688
rect 172334 131200 172390 131209
rect 172334 131135 172390 131144
rect 171322 130656 171378 130665
rect 171322 130591 171378 130600
rect 171336 126954 171364 130591
rect 172242 130112 172298 130121
rect 172242 130047 172298 130056
rect 172256 130014 172284 130047
rect 172244 130008 172296 130014
rect 172244 129950 172296 129956
rect 172150 129024 172206 129033
rect 172150 128959 172206 128968
rect 171966 128480 172022 128489
rect 171966 128415 172022 128424
rect 171782 127392 171838 127401
rect 171782 127327 171838 127336
rect 171324 126948 171376 126954
rect 171324 126890 171376 126896
rect 171506 125216 171562 125225
rect 171506 125151 171562 125160
rect 171520 124370 171548 125151
rect 171508 124364 171560 124370
rect 171508 124306 171560 124312
rect 170404 122800 170456 122806
rect 170404 122742 170456 122748
rect 171796 114510 171824 127327
rect 171874 124672 171930 124681
rect 171874 124607 171930 124616
rect 171888 124302 171916 124607
rect 171876 124296 171928 124302
rect 171876 124238 171928 124244
rect 171980 124114 172008 128415
rect 172058 127936 172114 127945
rect 172058 127871 172114 127880
rect 171888 124086 172008 124114
rect 171888 118658 171916 124086
rect 172072 123978 172100 127871
rect 172164 125610 172192 128959
rect 172348 128314 172376 131135
rect 172440 131102 172468 131679
rect 172428 131096 172480 131102
rect 172428 131038 172480 131044
rect 172426 129568 172482 129577
rect 172482 129526 172560 129554
rect 172426 129503 172482 129512
rect 172336 128308 172388 128314
rect 172336 128250 172388 128256
rect 172334 126848 172390 126857
rect 172334 126783 172390 126792
rect 172244 125792 172296 125798
rect 172242 125760 172244 125769
rect 172296 125760 172298 125769
rect 172242 125695 172298 125704
rect 172348 125662 172376 126783
rect 172426 126304 172482 126313
rect 172426 126239 172482 126248
rect 172440 125730 172468 126239
rect 172428 125724 172480 125730
rect 172428 125666 172480 125672
rect 172336 125656 172388 125662
rect 172164 125582 172284 125610
rect 172336 125598 172388 125604
rect 172150 124264 172206 124273
rect 172150 124199 172152 124208
rect 172204 124199 172206 124208
rect 172152 124170 172204 124176
rect 171980 123950 172100 123978
rect 171876 118652 171928 118658
rect 171876 118594 171928 118600
rect 171980 115938 172008 123950
rect 172256 122834 172284 125582
rect 172532 124914 172560 129526
rect 172520 124908 172572 124914
rect 172520 124850 172572 124856
rect 175924 124364 175976 124370
rect 175924 124306 175976 124312
rect 174544 124296 174596 124302
rect 174544 124238 174596 124244
rect 173164 124228 173216 124234
rect 173164 124170 173216 124176
rect 172072 122806 172284 122834
rect 172072 120086 172100 122806
rect 172060 120080 172112 120086
rect 172060 120022 172112 120028
rect 171968 115932 172020 115938
rect 171968 115874 172020 115880
rect 171784 114504 171836 114510
rect 171784 114446 171836 114452
rect 173176 102134 173204 124170
rect 174556 103494 174584 124238
rect 175936 112470 175964 124306
rect 177316 122942 177344 224946
rect 177408 172446 177436 247046
rect 177396 172440 177448 172446
rect 177396 172382 177448 172388
rect 178696 160750 178724 287030
rect 198186 286240 198242 286249
rect 198186 286175 198242 286184
rect 197358 284200 197414 284209
rect 197358 284135 197414 284144
rect 197372 282946 197400 284135
rect 197360 282940 197412 282946
rect 197360 282882 197412 282888
rect 197910 282024 197966 282033
rect 197910 281959 197966 281968
rect 197924 281586 197952 281959
rect 197912 281580 197964 281586
rect 197912 281522 197964 281528
rect 197542 279984 197598 279993
rect 197542 279919 197598 279928
rect 197556 278798 197584 279919
rect 197544 278792 197596 278798
rect 197544 278734 197596 278740
rect 197358 277808 197414 277817
rect 197358 277743 197414 277752
rect 197372 277438 197400 277743
rect 181444 277432 181496 277438
rect 181444 277374 181496 277380
rect 197360 277432 197412 277438
rect 197360 277374 197412 277380
rect 180064 273284 180116 273290
rect 180064 273226 180116 273232
rect 178776 258120 178828 258126
rect 178776 258062 178828 258068
rect 178788 177954 178816 258062
rect 180076 186250 180104 273226
rect 180156 260908 180208 260914
rect 180156 260850 180208 260856
rect 180064 186244 180116 186250
rect 180064 186186 180116 186192
rect 178868 182232 178920 182238
rect 178868 182174 178920 182180
rect 178776 177948 178828 177954
rect 178776 177890 178828 177896
rect 178776 167680 178828 167686
rect 178776 167622 178828 167628
rect 178684 160744 178736 160750
rect 178684 160686 178736 160692
rect 177396 158772 177448 158778
rect 177396 158714 177448 158720
rect 177408 139330 177436 158714
rect 178788 141982 178816 167622
rect 178880 145858 178908 182174
rect 180168 179246 180196 260850
rect 180248 205692 180300 205698
rect 180248 205634 180300 205640
rect 180156 179240 180208 179246
rect 180156 179182 180208 179188
rect 180064 162920 180116 162926
rect 180064 162862 180116 162868
rect 178868 145852 178920 145858
rect 178868 145794 178920 145800
rect 179420 142180 179472 142186
rect 179420 142122 179472 142128
rect 178776 141976 178828 141982
rect 178776 141918 178828 141924
rect 178040 140820 178092 140826
rect 178040 140762 178092 140768
rect 177396 139324 177448 139330
rect 177396 139266 177448 139272
rect 178052 135182 178080 140762
rect 179432 135318 179460 142122
rect 180076 141302 180104 162862
rect 180260 151502 180288 205634
rect 181456 189038 181484 277374
rect 197542 275768 197598 275777
rect 197542 275703 197598 275712
rect 197556 274718 197584 275703
rect 188344 274712 188396 274718
rect 188344 274654 188396 274660
rect 197544 274712 197596 274718
rect 197544 274654 197596 274660
rect 186964 270564 187016 270570
rect 186964 270506 187016 270512
rect 184204 266416 184256 266422
rect 184204 266358 184256 266364
rect 182824 264988 182876 264994
rect 182824 264930 182876 264936
rect 181536 262268 181588 262274
rect 181536 262210 181588 262216
rect 181444 189032 181496 189038
rect 181444 188974 181496 188980
rect 181548 180810 181576 262210
rect 181628 207052 181680 207058
rect 181628 206994 181680 207000
rect 181536 180804 181588 180810
rect 181536 180746 181588 180752
rect 180340 178084 180392 178090
rect 180340 178026 180392 178032
rect 180352 163674 180380 178026
rect 180340 163668 180392 163674
rect 180340 163610 180392 163616
rect 181444 162172 181496 162178
rect 181444 162114 181496 162120
rect 180248 151496 180300 151502
rect 180248 151438 180300 151444
rect 181456 142118 181484 162114
rect 181640 151774 181668 206994
rect 182836 182170 182864 264930
rect 182916 209840 182968 209846
rect 182916 209782 182968 209788
rect 182824 182164 182876 182170
rect 182824 182106 182876 182112
rect 182824 167068 182876 167074
rect 182824 167010 182876 167016
rect 181628 151768 181680 151774
rect 181628 151710 181680 151716
rect 181536 144968 181588 144974
rect 181536 144910 181588 144916
rect 181444 142112 181496 142118
rect 181444 142054 181496 142060
rect 180064 141296 180116 141302
rect 180064 141238 180116 141244
rect 181548 136542 181576 144910
rect 182836 142866 182864 167010
rect 182928 153134 182956 209782
rect 184216 183530 184244 266358
rect 184296 211200 184348 211206
rect 184296 211142 184348 211148
rect 184204 183524 184256 183530
rect 184204 183466 184256 183472
rect 184204 172576 184256 172582
rect 184204 172518 184256 172524
rect 182916 153128 182968 153134
rect 182916 153070 182968 153076
rect 182916 146328 182968 146334
rect 182916 146270 182968 146276
rect 182824 142860 182876 142866
rect 182824 142802 182876 142808
rect 182928 136610 182956 146270
rect 184216 144226 184244 172518
rect 184308 153202 184336 211142
rect 186976 184822 187004 270506
rect 187056 213988 187108 213994
rect 187056 213930 187108 213936
rect 186964 184816 187016 184822
rect 186964 184758 187016 184764
rect 186964 173936 187016 173942
rect 186964 173878 187016 173884
rect 184296 153196 184348 153202
rect 184296 153138 184348 153144
rect 184296 149116 184348 149122
rect 184296 149058 184348 149064
rect 184204 144220 184256 144226
rect 184204 144162 184256 144168
rect 184308 137290 184336 149058
rect 186976 143546 187004 173878
rect 187068 154494 187096 213930
rect 188356 187678 188384 274654
rect 197358 273592 197414 273601
rect 197358 273527 197414 273536
rect 197372 273290 197400 273527
rect 197360 273284 197412 273290
rect 197360 273226 197412 273232
rect 197542 271552 197598 271561
rect 197542 271487 197598 271496
rect 197556 270570 197584 271487
rect 197544 270564 197596 270570
rect 197544 270506 197596 270512
rect 193864 269340 193916 269346
rect 193864 269282 193916 269288
rect 192576 251252 192628 251258
rect 192576 251194 192628 251200
rect 191196 249824 191248 249830
rect 191196 249766 191248 249772
rect 191104 220924 191156 220930
rect 191104 220866 191156 220872
rect 188436 216708 188488 216714
rect 188436 216650 188488 216656
rect 188344 187672 188396 187678
rect 188344 187614 188396 187620
rect 188344 176724 188396 176730
rect 188344 176666 188396 176672
rect 188356 156670 188384 176666
rect 188344 156664 188396 156670
rect 188344 156606 188396 156612
rect 188448 154562 188476 216650
rect 188436 154556 188488 154562
rect 188436 154498 188488 154504
rect 187056 154488 187108 154494
rect 187056 154430 187108 154436
rect 188344 153264 188396 153270
rect 188344 153206 188396 153212
rect 187056 150476 187108 150482
rect 187056 150418 187108 150424
rect 186964 143540 187016 143546
rect 186964 143482 187016 143488
rect 187068 140078 187096 150418
rect 187056 140072 187108 140078
rect 187056 140014 187108 140020
rect 188356 137970 188384 153206
rect 188344 137964 188396 137970
rect 188344 137906 188396 137912
rect 184296 137284 184348 137290
rect 184296 137226 184348 137232
rect 182916 136604 182968 136610
rect 182916 136546 182968 136552
rect 181536 136536 181588 136542
rect 181536 136478 181588 136484
rect 179420 135312 179472 135318
rect 179420 135254 179472 135260
rect 178040 135176 178092 135182
rect 178040 135118 178092 135124
rect 178040 130008 178092 130014
rect 178040 129950 178092 129956
rect 178052 124166 178080 129950
rect 180064 125792 180116 125798
rect 180064 125734 180116 125740
rect 178040 124160 178092 124166
rect 178040 124102 178092 124108
rect 177304 122936 177356 122942
rect 177304 122878 177356 122884
rect 175924 112464 175976 112470
rect 175924 112406 175976 112412
rect 180076 107642 180104 125734
rect 181444 125724 181496 125730
rect 181444 125666 181496 125672
rect 181456 110430 181484 125666
rect 182824 125656 182876 125662
rect 182824 125598 182876 125604
rect 182836 111790 182864 125598
rect 191116 122806 191144 220866
rect 191208 173874 191236 249766
rect 192484 218068 192536 218074
rect 192484 218010 192536 218016
rect 191196 173868 191248 173874
rect 191196 173810 191248 173816
rect 192496 122874 192524 218010
rect 192588 175234 192616 251194
rect 193876 184890 193904 269282
rect 197634 267336 197690 267345
rect 197634 267271 197690 267280
rect 197648 266422 197676 267271
rect 197636 266416 197688 266422
rect 197636 266358 197688 266364
rect 197358 265160 197414 265169
rect 197358 265095 197414 265104
rect 197372 264994 197400 265095
rect 197360 264988 197412 264994
rect 197360 264930 197412 264936
rect 197358 263120 197414 263129
rect 197358 263055 197414 263064
rect 197372 262274 197400 263055
rect 197360 262268 197412 262274
rect 197360 262210 197412 262216
rect 197358 260944 197414 260953
rect 197358 260879 197360 260888
rect 197412 260879 197414 260888
rect 197360 260850 197412 260856
rect 197358 258904 197414 258913
rect 197358 258839 197414 258848
rect 197372 258126 197400 258839
rect 197360 258120 197412 258126
rect 197360 258062 197412 258068
rect 196624 256760 196676 256766
rect 196624 256702 196676 256708
rect 195244 253972 195296 253978
rect 195244 253914 195296 253920
rect 193956 190936 194008 190942
rect 193956 190878 194008 190884
rect 193864 184884 193916 184890
rect 193864 184826 193916 184832
rect 192576 175228 192628 175234
rect 192576 175170 192628 175176
rect 193968 147626 193996 190878
rect 195256 176662 195284 253914
rect 195336 241528 195388 241534
rect 195336 241470 195388 241476
rect 195244 176656 195296 176662
rect 195244 176598 195296 176604
rect 195348 169726 195376 241470
rect 195428 180940 195480 180946
rect 195428 180882 195480 180888
rect 195336 169720 195388 169726
rect 195336 169662 195388 169668
rect 193956 147620 194008 147626
rect 193956 147562 194008 147568
rect 195440 144906 195468 180882
rect 196636 178022 196664 256702
rect 198002 254688 198058 254697
rect 198002 254623 198058 254632
rect 198016 253978 198044 254623
rect 198004 253972 198056 253978
rect 198004 253914 198056 253920
rect 197910 252512 197966 252521
rect 197910 252447 197966 252456
rect 197924 251258 197952 252447
rect 197912 251252 197964 251258
rect 197912 251194 197964 251200
rect 198094 250472 198150 250481
rect 198094 250407 198150 250416
rect 198108 249830 198136 250407
rect 198096 249824 198148 249830
rect 198096 249766 198148 249772
rect 197542 248296 197598 248305
rect 197542 248231 197598 248240
rect 197556 247110 197584 248231
rect 197544 247104 197596 247110
rect 197544 247046 197596 247052
rect 198094 246256 198150 246265
rect 198094 246191 198150 246200
rect 197542 244080 197598 244089
rect 197542 244015 197598 244024
rect 197556 242962 197584 244015
rect 197544 242956 197596 242962
rect 197544 242898 197596 242904
rect 197542 239864 197598 239873
rect 197542 239799 197598 239808
rect 197556 238814 197584 239799
rect 197544 238808 197596 238814
rect 197544 238750 197596 238756
rect 196716 237788 196768 237794
rect 196716 237730 196768 237736
rect 196624 178016 196676 178022
rect 196624 177958 196676 177964
rect 196728 167006 196756 237730
rect 197542 235648 197598 235657
rect 197542 235583 197598 235592
rect 197556 234666 197584 235583
rect 197544 234660 197596 234666
rect 197544 234602 197596 234608
rect 197358 233608 197414 233617
rect 197358 233543 197414 233552
rect 197372 233306 197400 233543
rect 197360 233300 197412 233306
rect 197360 233242 197412 233248
rect 197358 229392 197414 229401
rect 197358 229327 197414 229336
rect 197372 229158 197400 229327
rect 197360 229152 197412 229158
rect 197360 229094 197412 229100
rect 197542 227352 197598 227361
rect 197542 227287 197598 227296
rect 197556 226370 197584 227287
rect 197544 226364 197596 226370
rect 197544 226306 197596 226312
rect 197358 225176 197414 225185
rect 197358 225111 197414 225120
rect 197372 225010 197400 225111
rect 197360 225004 197412 225010
rect 197360 224946 197412 224952
rect 198002 223136 198058 223145
rect 198002 223071 198058 223080
rect 197358 220960 197414 220969
rect 197358 220895 197360 220904
rect 197412 220895 197414 220904
rect 197360 220866 197412 220872
rect 197542 218920 197598 218929
rect 197542 218855 197598 218864
rect 197556 218074 197584 218855
rect 197544 218068 197596 218074
rect 197544 218010 197596 218016
rect 197358 216744 197414 216753
rect 197358 216679 197360 216688
rect 197412 216679 197414 216688
rect 197360 216650 197412 216656
rect 197358 214704 197414 214713
rect 197358 214639 197414 214648
rect 197372 213994 197400 214639
rect 197360 213988 197412 213994
rect 197360 213930 197412 213936
rect 197358 212528 197414 212537
rect 197358 212463 197414 212472
rect 197372 211206 197400 212463
rect 197360 211200 197412 211206
rect 197360 211142 197412 211148
rect 197358 210488 197414 210497
rect 197358 210423 197414 210432
rect 197372 209846 197400 210423
rect 197360 209840 197412 209846
rect 197360 209782 197412 209788
rect 197358 208312 197414 208321
rect 197358 208247 197414 208256
rect 197372 207058 197400 208247
rect 197360 207052 197412 207058
rect 197360 206994 197412 207000
rect 197358 206272 197414 206281
rect 197358 206207 197414 206216
rect 197372 205698 197400 206207
rect 197360 205692 197412 205698
rect 197360 205634 197412 205640
rect 197358 202056 197414 202065
rect 197358 201991 197414 202000
rect 197372 201550 197400 201991
rect 197360 201544 197412 201550
rect 197360 201486 197412 201492
rect 197542 199880 197598 199889
rect 197542 199815 197598 199824
rect 197556 198762 197584 199815
rect 197544 198756 197596 198762
rect 197544 198698 197596 198704
rect 197358 197840 197414 197849
rect 197358 197775 197414 197784
rect 197372 197402 197400 197775
rect 197360 197396 197412 197402
rect 197360 197338 197412 197344
rect 197542 195664 197598 195673
rect 197542 195599 197598 195608
rect 197556 194614 197584 195599
rect 197544 194608 197596 194614
rect 197544 194550 197596 194556
rect 197358 193624 197414 193633
rect 197358 193559 197414 193568
rect 197372 193254 197400 193559
rect 197360 193248 197412 193254
rect 197360 193190 197412 193196
rect 197358 189408 197414 189417
rect 197358 189343 197414 189352
rect 197372 189106 197400 189343
rect 197360 189100 197412 189106
rect 197360 189042 197412 189048
rect 197358 187232 197414 187241
rect 197358 187167 197414 187176
rect 197372 186386 197400 187167
rect 197360 186380 197412 186386
rect 197360 186322 197412 186328
rect 196808 185020 196860 185026
rect 196808 184962 196860 184968
rect 196716 167000 196768 167006
rect 196716 166942 196768 166948
rect 196820 146266 196848 184962
rect 197358 183016 197414 183025
rect 197358 182951 197414 182960
rect 197372 182238 197400 182951
rect 197360 182232 197412 182238
rect 197360 182174 197412 182180
rect 197358 178800 197414 178809
rect 197358 178735 197414 178744
rect 197372 178090 197400 178735
rect 197360 178084 197412 178090
rect 197360 178026 197412 178032
rect 197358 176760 197414 176769
rect 197358 176695 197360 176704
rect 197412 176695 197414 176704
rect 197360 176666 197412 176672
rect 197726 174584 197782 174593
rect 197726 174519 197782 174528
rect 197740 173942 197768 174519
rect 197728 173936 197780 173942
rect 197728 173878 197780 173884
rect 197360 172576 197412 172582
rect 197358 172544 197360 172553
rect 197412 172544 197414 172553
rect 197358 172479 197414 172488
rect 197450 170368 197506 170377
rect 197450 170303 197506 170312
rect 197358 168328 197414 168337
rect 197358 168263 197414 168272
rect 197372 167074 197400 168263
rect 197464 167686 197492 170303
rect 197452 167680 197504 167686
rect 197452 167622 197504 167628
rect 197360 167068 197412 167074
rect 197360 167010 197412 167016
rect 197542 164112 197598 164121
rect 197542 164047 197598 164056
rect 197556 162926 197584 164047
rect 197544 162920 197596 162926
rect 197544 162862 197596 162868
rect 197542 159896 197598 159905
rect 197542 159831 197598 159840
rect 197556 158778 197584 159831
rect 197544 158772 197596 158778
rect 197544 158714 197596 158720
rect 197358 157856 197414 157865
rect 197358 157791 197414 157800
rect 197372 157418 197400 157791
rect 197360 157412 197412 157418
rect 197360 157354 197412 157360
rect 197542 155680 197598 155689
rect 197542 155615 197598 155624
rect 197556 154630 197584 155615
rect 197544 154624 197596 154630
rect 197544 154566 197596 154572
rect 197358 153640 197414 153649
rect 197358 153575 197414 153584
rect 197372 153270 197400 153575
rect 197360 153264 197412 153270
rect 197360 153206 197412 153212
rect 197542 151464 197598 151473
rect 197542 151399 197598 151408
rect 197556 150482 197584 151399
rect 197544 150476 197596 150482
rect 197544 150418 197596 150424
rect 197358 149424 197414 149433
rect 197358 149359 197414 149368
rect 197372 149122 197400 149359
rect 197360 149116 197412 149122
rect 197360 149058 197412 149064
rect 197634 147248 197690 147257
rect 197634 147183 197690 147192
rect 197648 146334 197676 147183
rect 197636 146328 197688 146334
rect 197636 146270 197688 146276
rect 196808 146260 196860 146266
rect 196808 146202 196860 146208
rect 197358 145208 197414 145217
rect 197358 145143 197414 145152
rect 197372 144974 197400 145143
rect 197360 144968 197412 144974
rect 197360 144910 197412 144916
rect 195428 144900 195480 144906
rect 195428 144842 195480 144848
rect 197358 143032 197414 143041
rect 197358 142967 197414 142976
rect 197372 142186 197400 142967
rect 197360 142180 197412 142186
rect 197360 142122 197412 142128
rect 197358 140992 197414 141001
rect 197358 140927 197414 140936
rect 197372 140826 197400 140927
rect 197360 140820 197412 140826
rect 197360 140762 197412 140768
rect 197358 138816 197414 138825
rect 197358 138751 197414 138760
rect 197372 138038 197400 138751
rect 197360 138032 197412 138038
rect 197360 137974 197412 137980
rect 197358 136776 197414 136785
rect 197358 136711 197414 136720
rect 197372 136678 197400 136711
rect 197360 136672 197412 136678
rect 197360 136614 197412 136620
rect 198016 135930 198044 223071
rect 198108 171086 198136 246191
rect 198200 222902 198228 286175
rect 198462 269376 198518 269385
rect 198462 269311 198464 269320
rect 198516 269311 198518 269320
rect 198464 269282 198516 269288
rect 198372 256760 198424 256766
rect 198370 256728 198372 256737
rect 198424 256728 198426 256737
rect 198370 256663 198426 256672
rect 198278 242040 198334 242049
rect 198278 241975 198334 241984
rect 198292 241534 198320 241975
rect 198280 241528 198332 241534
rect 198280 241470 198332 241476
rect 198462 237824 198518 237833
rect 198462 237759 198464 237768
rect 198516 237759 198518 237768
rect 198464 237730 198516 237736
rect 198738 231568 198794 231577
rect 198738 231503 198794 231512
rect 198188 222896 198240 222902
rect 198188 222838 198240 222844
rect 198278 204096 198334 204105
rect 198278 204031 198334 204040
rect 198292 202910 198320 204031
rect 198280 202904 198332 202910
rect 198280 202846 198332 202852
rect 198278 191448 198334 191457
rect 198278 191383 198334 191392
rect 198292 190942 198320 191383
rect 198280 190936 198332 190942
rect 198280 190878 198332 190884
rect 198462 185192 198518 185201
rect 198462 185127 198518 185136
rect 198476 185026 198504 185127
rect 198464 185020 198516 185026
rect 198464 184962 198516 184968
rect 198278 180976 198334 180985
rect 198278 180911 198280 180920
rect 198332 180911 198334 180920
rect 198280 180882 198332 180888
rect 198096 171080 198148 171086
rect 198096 171022 198148 171028
rect 198462 166288 198518 166297
rect 198462 166223 198518 166232
rect 198476 162178 198504 166223
rect 198752 164218 198780 231503
rect 199396 215286 199424 301582
rect 201224 301368 201276 301374
rect 201224 301310 201276 301316
rect 200396 300892 200448 300898
rect 200396 300834 200448 300840
rect 200408 299948 200436 300834
rect 201236 299948 201264 301310
rect 202064 299948 202092 302398
rect 202880 300960 202932 300966
rect 202880 300902 202932 300908
rect 202892 299948 202920 300902
rect 203708 300144 203760 300150
rect 203708 300086 203760 300092
rect 203720 299948 203748 300086
rect 204640 299948 204668 303010
rect 206284 301436 206336 301442
rect 206284 301378 206336 301384
rect 205456 300212 205508 300218
rect 205456 300154 205508 300160
rect 205468 299948 205496 300154
rect 206296 299948 206324 301378
rect 207124 299948 207152 303078
rect 211344 302592 211396 302598
rect 211344 302534 211396 302540
rect 208860 302524 208912 302530
rect 208860 302466 208912 302472
rect 208872 299948 208900 302466
rect 210516 301572 210568 301578
rect 210516 301514 210568 301520
rect 210528 299948 210556 301514
rect 211356 299948 211384 302534
rect 212184 299948 212212 303146
rect 215576 301504 215628 301510
rect 215576 301446 215628 301452
rect 214748 301028 214800 301034
rect 214748 300970 214800 300976
rect 214760 299948 214788 300970
rect 215588 299948 215616 301446
rect 219360 299962 219388 324294
rect 220636 311908 220688 311914
rect 220636 311850 220688 311856
rect 220648 300286 220676 311850
rect 222120 306374 222148 378150
rect 221936 306346 222148 306374
rect 220728 304292 220780 304298
rect 220728 304234 220780 304240
rect 219808 300280 219860 300286
rect 219808 300222 219860 300228
rect 220636 300280 220688 300286
rect 220636 300222 220688 300228
rect 219006 299934 219388 299962
rect 219820 299948 219848 300222
rect 220740 299948 220768 304234
rect 221936 299962 221964 306346
rect 222384 304360 222436 304366
rect 222384 304302 222436 304308
rect 221582 299934 221964 299962
rect 222396 299948 222424 304302
rect 223408 299962 223436 404330
rect 224960 304496 225012 304502
rect 224960 304438 225012 304444
rect 224040 304428 224092 304434
rect 224040 304370 224092 304376
rect 223238 299934 223436 299962
rect 224052 299948 224080 304370
rect 224972 299948 225000 304438
rect 226168 299962 226196 456758
rect 226616 305652 226668 305658
rect 226616 305594 226668 305600
rect 225814 299934 226196 299962
rect 226628 299948 226656 305594
rect 227640 299962 227668 470562
rect 228272 305720 228324 305726
rect 228272 305662 228324 305668
rect 227470 299934 227668 299962
rect 228284 299948 228312 305662
rect 229192 302116 229244 302122
rect 229192 302058 229244 302064
rect 229204 299948 229232 302058
rect 230308 299962 230336 524418
rect 230400 302122 230428 536794
rect 230848 304564 230900 304570
rect 230848 304506 230900 304512
rect 230388 302116 230440 302122
rect 230388 302058 230440 302064
rect 230046 299934 230336 299962
rect 230860 299948 230888 304506
rect 231688 299948 231716 590650
rect 233160 304842 233188 699654
rect 237288 696992 237340 696998
rect 237288 696934 237340 696940
rect 235908 670744 235960 670750
rect 235908 670686 235960 670692
rect 234528 643136 234580 643142
rect 234528 643078 234580 643084
rect 234436 616888 234488 616894
rect 234436 616830 234488 616836
rect 233148 304836 233200 304842
rect 233148 304778 233200 304784
rect 232596 304632 232648 304638
rect 232596 304574 232648 304580
rect 232608 299948 232636 304574
rect 234448 300286 234476 616830
rect 233424 300280 233476 300286
rect 233424 300222 233476 300228
rect 234436 300280 234488 300286
rect 234436 300222 234488 300228
rect 233436 299948 233464 300222
rect 234540 299962 234568 643078
rect 235816 630692 235868 630698
rect 235816 630634 235868 630640
rect 235828 306374 235856 630634
rect 235552 306346 235856 306374
rect 235552 299962 235580 306346
rect 234278 299934 234568 299962
rect 235106 299934 235580 299962
rect 235920 299948 235948 670686
rect 237300 306374 237328 696934
rect 238576 683188 238628 683194
rect 238576 683130 238628 683136
rect 237208 306346 237328 306374
rect 237208 299962 237236 306346
rect 238484 304700 238536 304706
rect 238484 304642 238536 304648
rect 237656 300280 237708 300286
rect 237656 300222 237708 300228
rect 236854 299934 237236 299962
rect 237668 299948 237696 300222
rect 238496 299948 238524 304642
rect 238588 300286 238616 683130
rect 239312 307080 239364 307086
rect 239312 307022 239364 307028
rect 238576 300280 238628 300286
rect 238576 300222 238628 300228
rect 239324 299948 239352 307022
rect 241060 304768 241112 304774
rect 241060 304710 241112 304716
rect 240140 300280 240192 300286
rect 240140 300222 240192 300228
rect 240152 299948 240180 300222
rect 241072 299948 241100 304710
rect 241348 300286 241376 700266
rect 241888 307148 241940 307154
rect 241888 307090 241940 307096
rect 241336 300280 241388 300286
rect 241336 300222 241388 300228
rect 241900 299948 241928 307090
rect 242820 299962 242848 700470
rect 244464 307216 244516 307222
rect 244464 307158 244516 307164
rect 243544 305788 243596 305794
rect 243544 305730 243596 305736
rect 242742 299934 242848 299962
rect 243556 299948 243584 305730
rect 244476 299948 244504 307158
rect 245580 299962 245608 700674
rect 246948 330540 247000 330546
rect 246948 330482 247000 330488
rect 246120 305924 246172 305930
rect 246120 305866 246172 305872
rect 245318 299934 245608 299962
rect 246132 299948 246160 305866
rect 246960 299948 246988 330482
rect 248340 306374 248368 700878
rect 251088 700188 251140 700194
rect 251088 700130 251140 700136
rect 249708 700120 249760 700126
rect 249708 700062 249760 700068
rect 248248 306346 248368 306374
rect 248248 299962 248276 306346
rect 248696 306060 248748 306066
rect 248696 306002 248748 306008
rect 247802 299934 248276 299962
rect 248708 299948 248736 306002
rect 249720 299962 249748 700062
rect 251100 306374 251128 700130
rect 251192 325694 251220 700946
rect 255320 700868 255372 700874
rect 255320 700810 255372 700816
rect 253940 700800 253992 700806
rect 253940 700742 253992 700748
rect 252560 700256 252612 700262
rect 252560 700198 252612 700204
rect 251192 325666 251680 325694
rect 250824 306346 251128 306374
rect 250824 299962 250852 306346
rect 251180 304836 251232 304842
rect 251180 304778 251232 304784
rect 249550 299934 249748 299962
rect 250378 299934 250852 299962
rect 251192 299948 251220 304778
rect 251652 299962 251680 325666
rect 252572 299962 252600 700198
rect 253952 325694 253980 700742
rect 253952 325666 254256 325694
rect 253756 305992 253808 305998
rect 253756 305934 253808 305940
rect 251652 299934 252034 299962
rect 252572 299934 252954 299962
rect 253768 299948 253796 305934
rect 254228 299962 254256 325666
rect 255332 299962 255360 700810
rect 256792 700664 256844 700670
rect 256792 700606 256844 700612
rect 256700 700596 256752 700602
rect 256700 700538 256752 700544
rect 256712 306374 256740 700538
rect 256804 325694 256832 700606
rect 259552 700460 259604 700466
rect 259552 700402 259604 700408
rect 259460 700392 259512 700398
rect 259460 700334 259512 700340
rect 258080 327752 258132 327758
rect 258080 327694 258132 327700
rect 258092 325694 258120 327694
rect 256804 325666 257568 325694
rect 258092 325666 258488 325694
rect 256712 306346 256832 306374
rect 256240 305856 256292 305862
rect 256240 305798 256292 305804
rect 254228 299934 254610 299962
rect 255332 299934 255438 299962
rect 256252 299948 256280 305798
rect 256804 299962 256832 306346
rect 257540 299962 257568 325666
rect 258460 299962 258488 325666
rect 259472 299962 259500 700334
rect 259564 325694 259592 700402
rect 267660 700126 267688 703520
rect 283852 700194 283880 703520
rect 300136 700398 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 295984 700392 296036 700398
rect 295984 700334 296036 700340
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 283840 700188 283892 700194
rect 283840 700130 283892 700136
rect 267648 700120 267700 700126
rect 267648 700062 267700 700068
rect 260840 683256 260892 683262
rect 260840 683198 260892 683204
rect 260852 325694 260880 683198
rect 262220 670812 262272 670818
rect 262220 670754 262272 670760
rect 259564 325666 260144 325694
rect 260852 325666 261064 325694
rect 260116 299962 260144 325666
rect 261036 299962 261064 325666
rect 262232 303278 262260 670754
rect 262312 656940 262364 656946
rect 262312 656882 262364 656888
rect 262220 303272 262272 303278
rect 262220 303214 262272 303220
rect 262324 299962 262352 656882
rect 263600 632120 263652 632126
rect 263600 632062 263652 632068
rect 262772 303272 262824 303278
rect 262772 303214 262824 303220
rect 256804 299934 257186 299962
rect 257540 299934 258014 299962
rect 258460 299934 258842 299962
rect 259472 299934 259670 299962
rect 260116 299934 260590 299962
rect 261036 299934 261418 299962
rect 262246 299934 262352 299962
rect 262784 299962 262812 303214
rect 263612 299962 263640 632062
rect 264980 618316 265032 618322
rect 264980 618258 265032 618264
rect 263692 605872 263744 605878
rect 263692 605814 263744 605820
rect 263704 325694 263732 605814
rect 264992 325694 265020 618258
rect 266360 579692 266412 579698
rect 266360 579634 266412 579640
rect 263704 325666 264376 325694
rect 264992 325666 265296 325694
rect 264348 299962 264376 325666
rect 265268 299962 265296 325666
rect 266372 299962 266400 579634
rect 267740 565888 267792 565894
rect 267740 565830 267792 565836
rect 266452 553444 266504 553450
rect 266452 553386 266504 553392
rect 266464 325694 266492 553386
rect 266464 325666 266952 325694
rect 266924 299962 266952 325666
rect 267752 299962 267780 565830
rect 267832 527196 267884 527202
rect 267832 527138 267884 527144
rect 267844 325694 267872 527138
rect 270500 514820 270552 514826
rect 270500 514762 270552 514768
rect 269120 501016 269172 501022
rect 269120 500958 269172 500964
rect 269132 325694 269160 500958
rect 267844 325666 268608 325694
rect 269132 325666 269528 325694
rect 268580 299962 268608 325666
rect 269500 299962 269528 325666
rect 270512 299962 270540 514762
rect 270592 474768 270644 474774
rect 270592 474710 270644 474716
rect 270604 325694 270632 474710
rect 273260 462392 273312 462398
rect 273260 462334 273312 462340
rect 271880 448588 271932 448594
rect 271880 448530 271932 448536
rect 271892 325694 271920 448530
rect 270604 325666 271184 325694
rect 271892 325666 272104 325694
rect 271156 299962 271184 325666
rect 272076 299962 272104 325666
rect 262784 299934 263074 299962
rect 263612 299934 263902 299962
rect 264348 299934 264822 299962
rect 265268 299934 265650 299962
rect 266372 299934 266478 299962
rect 266924 299934 267306 299962
rect 267752 299934 268134 299962
rect 268580 299934 269054 299962
rect 269500 299934 269882 299962
rect 270512 299934 270710 299962
rect 271156 299934 271538 299962
rect 272076 299934 272458 299962
rect 273272 299948 273300 462334
rect 273352 422340 273404 422346
rect 273352 422282 273404 422288
rect 273364 325694 273392 422282
rect 274640 409896 274692 409902
rect 274640 409838 274692 409844
rect 273364 325666 273760 325694
rect 273732 299962 273760 325666
rect 274652 303278 274680 409838
rect 274732 397520 274784 397526
rect 274732 397462 274784 397468
rect 274640 303272 274692 303278
rect 274640 303214 274692 303220
rect 274744 299962 274772 397462
rect 276020 371272 276072 371278
rect 276020 371214 276072 371220
rect 276032 325694 276060 371214
rect 277400 357468 277452 357474
rect 277400 357410 277452 357416
rect 276032 325666 276336 325694
rect 275468 303272 275520 303278
rect 275468 303214 275520 303220
rect 275480 299962 275508 303214
rect 276308 299962 276336 325666
rect 277412 303278 277440 357410
rect 277492 345092 277544 345098
rect 277492 345034 277544 345040
rect 277400 303272 277452 303278
rect 277400 303214 277452 303220
rect 273732 299934 274114 299962
rect 274744 299934 274942 299962
rect 275480 299934 275770 299962
rect 276308 299934 276690 299962
rect 277504 299948 277532 345034
rect 278780 318844 278832 318850
rect 278780 318786 278832 318792
rect 278044 303272 278096 303278
rect 278044 303214 278096 303220
rect 278056 299962 278084 303214
rect 278792 299962 278820 318786
rect 295996 306066 296024 700334
rect 302884 554124 302936 554130
rect 302884 554066 302936 554072
rect 300768 337408 300820 337414
rect 300768 337350 300820 337356
rect 295984 306060 296036 306066
rect 295984 306002 296036 306008
rect 280896 305040 280948 305046
rect 280896 304982 280948 304988
rect 278056 299934 278346 299962
rect 278792 299934 279174 299962
rect 280908 299948 280936 304982
rect 296076 303000 296128 303006
rect 296076 302942 296128 302948
rect 285956 302932 286008 302938
rect 285956 302874 286008 302880
rect 284208 301640 284260 301646
rect 284208 301582 284260 301588
rect 281724 301096 281776 301102
rect 281724 301038 281776 301044
rect 281736 299948 281764 301038
rect 284220 299948 284248 301582
rect 284852 300076 284904 300082
rect 284852 300018 284904 300024
rect 284864 299962 284892 300018
rect 284864 299934 285154 299962
rect 285968 299948 285996 302874
rect 288532 302864 288584 302870
rect 288532 302806 288584 302812
rect 287612 301300 287664 301306
rect 287612 301242 287664 301248
rect 287624 299948 287652 301242
rect 288544 299948 288572 302806
rect 293592 302796 293644 302802
rect 293592 302738 293644 302744
rect 291016 302660 291068 302666
rect 291016 302602 291068 302608
rect 289084 300008 289136 300014
rect 289136 299956 289386 299962
rect 289084 299950 289386 299956
rect 289096 299934 289386 299950
rect 291028 299948 291056 302602
rect 292764 301164 292816 301170
rect 292764 301106 292816 301112
rect 291488 299946 291870 299962
rect 292776 299948 292804 301106
rect 293604 299948 293632 302738
rect 295248 302728 295300 302734
rect 295248 302670 295300 302676
rect 294420 301232 294472 301238
rect 294420 301174 294472 301180
rect 294432 299948 294460 301174
rect 295260 299948 295288 302670
rect 296088 299948 296116 302942
rect 300780 302870 300808 337350
rect 299480 302864 299532 302870
rect 299480 302806 299532 302812
rect 300768 302864 300820 302870
rect 300768 302806 300820 302812
rect 296996 302388 297048 302394
rect 296996 302330 297048 302336
rect 297008 299948 297036 302330
rect 297824 302320 297876 302326
rect 297824 302262 297876 302268
rect 297836 299948 297864 302262
rect 298652 302252 298704 302258
rect 298652 302194 298704 302200
rect 298664 299948 298692 302194
rect 299492 299948 299520 302806
rect 301504 301572 301556 301578
rect 301504 301514 301556 301520
rect 291476 299940 291870 299946
rect 291528 299934 291870 299940
rect 291476 299882 291528 299888
rect 289820 299872 289872 299878
rect 286520 299810 286810 299826
rect 289872 299820 290214 299826
rect 289820 299814 290214 299820
rect 286508 299804 286810 299810
rect 286560 299798 286810 299804
rect 289832 299798 290214 299814
rect 286508 299746 286560 299752
rect 213368 299736 213420 299742
rect 209714 299674 210096 299690
rect 213118 299684 213368 299690
rect 213118 299678 213420 299684
rect 209714 299668 210108 299674
rect 209714 299662 210056 299668
rect 213118 299662 213408 299678
rect 210056 299610 210108 299616
rect 208216 299600 208268 299606
rect 207966 299548 208216 299554
rect 207966 299542 208268 299548
rect 207966 299526 208256 299542
rect 218178 299538 218560 299554
rect 218178 299532 218572 299538
rect 218178 299526 218520 299532
rect 218520 299474 218572 299480
rect 214012 299464 214064 299470
rect 213826 299432 213882 299441
rect 213882 299390 213946 299418
rect 282644 299464 282696 299470
rect 216034 299432 216090 299441
rect 214012 299406 214064 299412
rect 213826 299367 213882 299376
rect 214024 299334 214052 299406
rect 214484 299390 214696 299418
rect 214012 299328 214064 299334
rect 214012 299270 214064 299276
rect 214378 299296 214434 299305
rect 214484 299282 214512 299390
rect 214668 299334 214696 299390
rect 216034 299367 216090 299376
rect 216954 299432 217010 299441
rect 282644 299406 282696 299412
rect 283472 299464 283524 299470
rect 283472 299406 283524 299412
rect 216954 299367 217010 299376
rect 216048 299334 216076 299367
rect 216968 299334 216996 299367
rect 282656 299334 282684 299406
rect 283484 299334 283512 299406
rect 214564 299328 214616 299334
rect 214434 299254 214512 299282
rect 214562 299296 214564 299305
rect 214656 299328 214708 299334
rect 214616 299296 214618 299305
rect 214378 299231 214434 299240
rect 214656 299270 214708 299276
rect 216036 299328 216088 299334
rect 216864 299328 216916 299334
rect 216036 299270 216088 299276
rect 216522 299276 216864 299282
rect 216522 299270 216916 299276
rect 216956 299328 217008 299334
rect 217600 299328 217652 299334
rect 216956 299270 217008 299276
rect 217350 299276 217600 299282
rect 224408 299328 224460 299334
rect 217350 299270 217652 299276
rect 224406 299296 224408 299305
rect 279700 299328 279752 299334
rect 224460 299296 224462 299305
rect 216522 299254 216904 299270
rect 217350 299254 217640 299270
rect 214562 299231 214618 299240
rect 282276 299328 282328 299334
rect 279752 299276 280002 299282
rect 279700 299270 280002 299276
rect 282644 299328 282696 299334
rect 282328 299276 282578 299282
rect 282276 299270 282578 299276
rect 282644 299270 282696 299276
rect 283012 299328 283064 299334
rect 283472 299328 283524 299334
rect 283064 299276 283406 299282
rect 283012 299270 283406 299276
rect 283472 299270 283524 299276
rect 279712 299254 280002 299270
rect 282288 299254 282578 299270
rect 283024 299254 283406 299270
rect 224406 299231 224462 299240
rect 199384 215280 199436 215286
rect 199384 215222 199436 215228
rect 301516 167006 301544 301514
rect 302896 298489 302924 554066
rect 323584 482452 323636 482458
rect 323584 482394 323636 482400
rect 302976 482384 303028 482390
rect 302976 482326 303028 482332
rect 302882 298480 302938 298489
rect 302882 298415 302938 298424
rect 302884 297424 302936 297430
rect 302884 297366 302936 297372
rect 302792 295384 302844 295390
rect 302790 295352 302792 295361
rect 302844 295352 302846 295361
rect 302790 295287 302846 295296
rect 302240 289264 302292 289270
rect 302238 289232 302240 289241
rect 302292 289232 302294 289241
rect 302238 289167 302294 289176
rect 302240 286544 302292 286550
rect 302240 286486 302292 286492
rect 302252 286113 302280 286486
rect 302238 286104 302294 286113
rect 302238 286039 302294 286048
rect 302790 283112 302846 283121
rect 302790 283047 302846 283056
rect 302804 282946 302832 283047
rect 302792 282940 302844 282946
rect 302792 282882 302844 282888
rect 302422 279984 302478 279993
rect 302422 279919 302478 279928
rect 302436 278798 302464 279919
rect 302424 278792 302476 278798
rect 302424 278734 302476 278740
rect 302790 276856 302846 276865
rect 302790 276791 302846 276800
rect 302804 276078 302832 276791
rect 302792 276072 302844 276078
rect 302792 276014 302844 276020
rect 302698 273864 302754 273873
rect 302698 273799 302754 273808
rect 302712 273290 302740 273799
rect 302700 273284 302752 273290
rect 302700 273226 302752 273232
rect 302896 267753 302924 297366
rect 302988 292369 303016 482326
rect 304264 409216 304316 409222
rect 304264 409158 304316 409164
rect 303068 297492 303120 297498
rect 303068 297434 303120 297440
rect 302974 292360 303030 292369
rect 302974 292295 303030 292304
rect 303080 270745 303108 297434
rect 304276 286550 304304 409158
rect 304356 409148 304408 409154
rect 304356 409090 304408 409096
rect 304368 289270 304396 409090
rect 322204 337476 322256 337482
rect 322204 337418 322256 337424
rect 307024 302320 307076 302326
rect 307024 302262 307076 302268
rect 305644 302252 305696 302258
rect 305644 302194 305696 302200
rect 304356 289264 304408 289270
rect 304356 289206 304408 289212
rect 304264 286544 304316 286550
rect 304264 286486 304316 286492
rect 303066 270736 303122 270745
rect 303066 270671 303122 270680
rect 303344 268456 303396 268462
rect 303344 268398 303396 268404
rect 303252 268388 303304 268394
rect 303252 268330 303304 268336
rect 302882 267744 302938 267753
rect 302882 267679 302938 267688
rect 303160 267028 303212 267034
rect 303160 266970 303212 266976
rect 302700 264920 302752 264926
rect 302700 264862 302752 264868
rect 302712 264625 302740 264862
rect 302698 264616 302754 264625
rect 302698 264551 302754 264560
rect 302884 264240 302936 264246
rect 302884 264182 302936 264188
rect 302332 262200 302384 262206
rect 302332 262142 302384 262148
rect 302344 261497 302372 262142
rect 302330 261488 302386 261497
rect 302330 261423 302386 261432
rect 302606 258496 302662 258505
rect 302606 258431 302662 258440
rect 302620 258126 302648 258431
rect 302608 258120 302660 258126
rect 302608 258062 302660 258068
rect 302792 256012 302844 256018
rect 302792 255954 302844 255960
rect 302804 255377 302832 255954
rect 302790 255368 302846 255377
rect 302790 255303 302846 255312
rect 302790 249248 302846 249257
rect 302790 249183 302846 249192
rect 302804 248470 302832 249183
rect 302792 248464 302844 248470
rect 302792 248406 302844 248412
rect 302514 246120 302570 246129
rect 302514 246055 302570 246064
rect 302528 245682 302556 246055
rect 302516 245676 302568 245682
rect 302516 245618 302568 245624
rect 302896 240009 302924 264182
rect 303172 258074 303200 266970
rect 303264 265010 303292 268330
rect 303356 267734 303384 268398
rect 303356 267706 303568 267734
rect 303264 264982 303384 265010
rect 303172 258046 303292 258074
rect 303264 252249 303292 258046
rect 302974 252240 303030 252249
rect 302974 252175 303030 252184
rect 303250 252240 303306 252249
rect 303250 252175 303306 252184
rect 302988 251258 303016 252175
rect 302976 251252 303028 251258
rect 302976 251194 303028 251200
rect 303356 251138 303384 264982
rect 303264 251110 303384 251138
rect 303264 243137 303292 251110
rect 303344 250504 303396 250510
rect 303344 250446 303396 250452
rect 303356 248414 303384 250446
rect 303356 248386 303476 248414
rect 303250 243128 303306 243137
rect 303250 243063 303306 243072
rect 303264 242962 303292 243063
rect 303252 242956 303304 242962
rect 303252 242898 303304 242904
rect 302882 240000 302938 240009
rect 302882 239935 302938 239944
rect 302790 236872 302846 236881
rect 302790 236807 302846 236816
rect 302804 236026 302832 236807
rect 302792 236020 302844 236026
rect 302792 235962 302844 235968
rect 302698 233880 302754 233889
rect 302698 233815 302754 233824
rect 302712 233306 302740 233815
rect 302700 233300 302752 233306
rect 302700 233242 302752 233248
rect 302790 230752 302846 230761
rect 302790 230687 302846 230696
rect 302804 230518 302832 230687
rect 302792 230512 302844 230518
rect 302792 230454 302844 230460
rect 302792 227724 302844 227730
rect 302792 227666 302844 227672
rect 302804 227633 302832 227666
rect 302790 227624 302846 227633
rect 302790 227559 302846 227568
rect 302330 224632 302386 224641
rect 302330 224567 302386 224576
rect 302344 223990 302372 224567
rect 302896 224398 302924 239935
rect 303264 238754 303292 242898
rect 303264 238726 303384 238754
rect 302976 225616 303028 225622
rect 302976 225558 303028 225564
rect 302884 224392 302936 224398
rect 302884 224334 302936 224340
rect 302884 224256 302936 224262
rect 302884 224198 302936 224204
rect 302332 223984 302384 223990
rect 302332 223926 302384 223932
rect 302332 222148 302384 222154
rect 302332 222090 302384 222096
rect 302344 221513 302372 222090
rect 302330 221504 302386 221513
rect 302330 221439 302386 221448
rect 302424 219428 302476 219434
rect 302424 219370 302476 219376
rect 302436 218385 302464 219370
rect 302422 218376 302478 218385
rect 302422 218311 302478 218320
rect 302896 212265 302924 224198
rect 302882 212256 302938 212265
rect 302882 212191 302938 212200
rect 302240 206168 302292 206174
rect 302238 206136 302240 206145
rect 302292 206136 302294 206145
rect 302238 206071 302294 206080
rect 302790 196888 302846 196897
rect 302790 196823 302846 196832
rect 302804 196654 302832 196823
rect 302792 196648 302844 196654
rect 302792 196590 302844 196596
rect 302606 193760 302662 193769
rect 302606 193695 302662 193704
rect 302620 193254 302648 193695
rect 302608 193248 302660 193254
rect 302608 193190 302660 193196
rect 302424 191820 302476 191826
rect 302424 191762 302476 191768
rect 302436 190777 302464 191762
rect 302422 190768 302478 190777
rect 302422 190703 302478 190712
rect 302792 184884 302844 184890
rect 302792 184826 302844 184832
rect 302804 184657 302832 184826
rect 302790 184648 302846 184657
rect 302790 184583 302846 184592
rect 302700 182164 302752 182170
rect 302700 182106 302752 182112
rect 302712 181529 302740 182106
rect 302698 181520 302754 181529
rect 302698 181455 302754 181464
rect 302238 175400 302294 175409
rect 302238 175335 302294 175344
rect 302252 175302 302280 175335
rect 302240 175296 302292 175302
rect 302240 175238 302292 175244
rect 302790 169144 302846 169153
rect 302790 169079 302846 169088
rect 302804 169046 302832 169079
rect 302792 169040 302844 169046
rect 302792 168982 302844 168988
rect 301504 167000 301556 167006
rect 301504 166942 301556 166948
rect 302792 166320 302844 166326
rect 302792 166262 302844 166268
rect 302804 166161 302832 166262
rect 302790 166152 302846 166161
rect 302790 166087 302846 166096
rect 198740 164212 198792 164218
rect 198740 164154 198792 164160
rect 302790 163024 302846 163033
rect 302790 162959 302846 162968
rect 302804 162926 302832 162959
rect 302792 162920 302844 162926
rect 302792 162862 302844 162868
rect 198464 162172 198516 162178
rect 198464 162114 198516 162120
rect 198094 162072 198150 162081
rect 198094 162007 198150 162016
rect 198108 148374 198136 162007
rect 302514 159896 302570 159905
rect 302514 159831 302570 159840
rect 302528 158778 302556 159831
rect 302516 158772 302568 158778
rect 302516 158714 302568 158720
rect 302896 158030 302924 212191
rect 302988 203017 303016 225558
rect 303068 215960 303120 215966
rect 303068 215902 303120 215908
rect 303080 215393 303108 215902
rect 303066 215384 303122 215393
rect 303066 215319 303122 215328
rect 303066 209264 303122 209273
rect 303066 209199 303122 209208
rect 303080 209098 303108 209199
rect 303068 209092 303120 209098
rect 303068 209034 303120 209040
rect 302974 203008 303030 203017
rect 302974 202943 303030 202952
rect 302884 158024 302936 158030
rect 302884 157966 302936 157972
rect 302790 156904 302846 156913
rect 302790 156839 302846 156848
rect 302804 153950 302832 156839
rect 302988 155242 303016 202943
rect 303356 195294 303384 238726
rect 303448 200025 303476 248386
rect 303540 215966 303568 267706
rect 304264 240780 304316 240786
rect 304264 240722 304316 240728
rect 303528 215960 303580 215966
rect 303528 215902 303580 215908
rect 303528 209092 303580 209098
rect 303528 209034 303580 209040
rect 303434 200016 303490 200025
rect 303434 199951 303490 199960
rect 303448 199442 303476 199951
rect 303436 199436 303488 199442
rect 303436 199378 303488 199384
rect 303344 195288 303396 195294
rect 303344 195230 303396 195236
rect 303066 187640 303122 187649
rect 303066 187575 303122 187584
rect 303080 186998 303108 187575
rect 303068 186992 303120 186998
rect 303068 186934 303120 186940
rect 303436 186992 303488 186998
rect 303436 186934 303488 186940
rect 303344 179376 303396 179382
rect 303344 179318 303396 179324
rect 303356 178401 303384 179318
rect 303342 178392 303398 178401
rect 303342 178327 303398 178336
rect 303066 172272 303122 172281
rect 303066 172207 303122 172216
rect 302976 155236 303028 155242
rect 302976 155178 303028 155184
rect 302792 153944 302844 153950
rect 302792 153886 302844 153892
rect 302790 153776 302846 153785
rect 302790 153711 302846 153720
rect 302700 153264 302752 153270
rect 302700 153206 302752 153212
rect 198096 148368 198148 148374
rect 198096 148310 198148 148316
rect 302712 147665 302740 153206
rect 302804 152590 302832 153711
rect 303080 152658 303108 172207
rect 303068 152652 303120 152658
rect 303068 152594 303120 152600
rect 302792 152584 302844 152590
rect 302792 152526 302844 152532
rect 303448 152522 303476 186934
rect 303540 153882 303568 209034
rect 304276 206174 304304 240722
rect 304908 225684 304960 225690
rect 304908 225626 304960 225632
rect 304264 206168 304316 206174
rect 304264 206110 304316 206116
rect 304920 179382 304948 225626
rect 305656 194546 305684 302194
rect 307036 266150 307064 302262
rect 309784 302252 309836 302258
rect 309784 302194 309836 302200
rect 307024 266144 307076 266150
rect 307024 266086 307076 266092
rect 307668 251252 307720 251258
rect 307668 251194 307720 251200
rect 305644 194540 305696 194546
rect 305644 194482 305696 194488
rect 305736 193860 305788 193866
rect 305736 193802 305788 193808
rect 304908 179376 304960 179382
rect 304908 179318 304960 179324
rect 303528 153876 303580 153882
rect 303528 153818 303580 153824
rect 303436 152516 303488 152522
rect 303436 152458 303488 152464
rect 302792 151768 302844 151774
rect 302792 151710 302844 151716
rect 302804 150793 302832 151710
rect 302790 150784 302846 150793
rect 302790 150719 302846 150728
rect 302698 147656 302754 147665
rect 302698 147591 302754 147600
rect 302792 144900 302844 144906
rect 302792 144842 302844 144848
rect 302804 144537 302832 144842
rect 302790 144528 302846 144537
rect 302790 144463 302846 144472
rect 302332 142112 302384 142118
rect 302332 142054 302384 142060
rect 302344 141545 302372 142054
rect 302330 141536 302386 141545
rect 302330 141471 302386 141480
rect 302882 138408 302938 138417
rect 302882 138343 302938 138352
rect 198004 135924 198056 135930
rect 198004 135866 198056 135872
rect 197726 134600 197782 134609
rect 197726 134535 197782 134544
rect 197740 133958 197768 134535
rect 197728 133952 197780 133958
rect 197728 133894 197780 133900
rect 197358 132560 197414 132569
rect 197358 132495 197360 132504
rect 197412 132495 197414 132504
rect 197360 132466 197412 132472
rect 302514 132288 302570 132297
rect 302514 132223 302570 132232
rect 197360 131096 197412 131102
rect 197360 131038 197412 131044
rect 197372 130393 197400 131038
rect 197358 130384 197414 130393
rect 197358 130319 197414 130328
rect 197358 128344 197414 128353
rect 197358 128279 197360 128288
rect 197412 128279 197414 128288
rect 197360 128250 197412 128256
rect 197636 126948 197688 126954
rect 197636 126890 197688 126896
rect 197648 126177 197676 126890
rect 197634 126168 197690 126177
rect 197634 126103 197690 126112
rect 302422 126168 302478 126177
rect 302422 126103 302478 126112
rect 302436 125254 302464 126103
rect 302424 125248 302476 125254
rect 302424 125190 302476 125196
rect 302528 125186 302556 132223
rect 302698 129160 302754 129169
rect 302698 129095 302754 129104
rect 302516 125180 302568 125186
rect 302516 125122 302568 125128
rect 302712 125050 302740 129095
rect 302896 125118 302924 138343
rect 302974 135280 303030 135289
rect 302974 135215 303030 135224
rect 302884 125112 302936 125118
rect 302884 125054 302936 125060
rect 302700 125044 302752 125050
rect 302700 124986 302752 124992
rect 302988 124982 303016 135215
rect 302976 124976 303028 124982
rect 302976 124918 303028 124924
rect 197452 124908 197504 124914
rect 197452 124850 197504 124856
rect 302240 124908 302292 124914
rect 302240 124850 302292 124856
rect 197360 124160 197412 124166
rect 197358 124128 197360 124137
rect 197412 124128 197414 124137
rect 197358 124063 197414 124072
rect 192484 122868 192536 122874
rect 192484 122810 192536 122816
rect 191104 122800 191156 122806
rect 191104 122742 191156 122748
rect 197464 121961 197492 124850
rect 302252 123049 302280 124850
rect 302976 123548 303028 123554
rect 302976 123490 303028 123496
rect 302884 123480 302936 123486
rect 302884 123422 302936 123428
rect 302238 123040 302294 123049
rect 302238 122975 302294 122984
rect 301504 122120 301556 122126
rect 301504 122062 301556 122068
rect 197450 121952 197506 121961
rect 197450 121887 197506 121896
rect 197360 120080 197412 120086
rect 197360 120022 197412 120028
rect 197372 119921 197400 120022
rect 197358 119912 197414 119921
rect 197358 119847 197414 119856
rect 197636 118652 197688 118658
rect 197636 118594 197688 118600
rect 197648 117745 197676 118594
rect 197634 117736 197690 117745
rect 197634 117671 197690 117680
rect 198556 115932 198608 115938
rect 198556 115874 198608 115880
rect 198568 115705 198596 115874
rect 198554 115696 198610 115705
rect 198554 115631 198610 115640
rect 197544 114504 197596 114510
rect 197544 114446 197596 114452
rect 197556 113529 197584 114446
rect 197542 113520 197598 113529
rect 197542 113455 197598 113464
rect 197452 112464 197504 112470
rect 197452 112406 197504 112412
rect 182824 111784 182876 111790
rect 182824 111726 182876 111732
rect 197360 111784 197412 111790
rect 197360 111726 197412 111732
rect 197372 111489 197400 111726
rect 197358 111480 197414 111489
rect 197358 111415 197414 111424
rect 181444 110424 181496 110430
rect 181444 110366 181496 110372
rect 180064 107636 180116 107642
rect 180064 107578 180116 107584
rect 197464 105097 197492 112406
rect 197544 110424 197596 110430
rect 197544 110366 197596 110372
rect 197556 109313 197584 110366
rect 197542 109304 197598 109313
rect 197542 109239 197598 109248
rect 198004 107636 198056 107642
rect 198004 107578 198056 107584
rect 198016 107273 198044 107578
rect 198002 107264 198058 107273
rect 198002 107199 198058 107208
rect 197450 105088 197506 105097
rect 197450 105023 197506 105032
rect 174544 103488 174596 103494
rect 174544 103430 174596 103436
rect 198004 103488 198056 103494
rect 198004 103430 198056 103436
rect 198016 103057 198044 103430
rect 198002 103048 198058 103057
rect 198002 102983 198058 102992
rect 173164 102128 173216 102134
rect 173164 102070 173216 102076
rect 198004 102128 198056 102134
rect 198004 102070 198056 102076
rect 198016 101017 198044 102070
rect 198002 101008 198058 101017
rect 198002 100943 198058 100952
rect 166908 99408 166960 99414
rect 166908 99350 166960 99356
rect 195334 97880 195390 97889
rect 195334 97815 195390 97824
rect 192484 97096 192536 97102
rect 192484 97038 192536 97044
rect 186964 96620 187016 96626
rect 186964 96562 187016 96568
rect 161388 96552 161440 96558
rect 161388 96494 161440 96500
rect 158628 95124 158680 95130
rect 158628 95066 158680 95072
rect 157984 71732 158036 71738
rect 157984 71674 158036 71680
rect 158640 3602 158668 95066
rect 160008 93832 160060 93838
rect 160008 93774 160060 93780
rect 160020 3602 160048 93774
rect 161204 14476 161256 14482
rect 161204 14418 161256 14424
rect 161216 3602 161244 14418
rect 161400 6914 161428 96494
rect 183468 96484 183520 96490
rect 183468 96426 183520 96432
rect 179328 96416 179380 96422
rect 179328 96358 179380 96364
rect 176568 96348 176620 96354
rect 176568 96290 176620 96296
rect 173164 96280 173216 96286
rect 173164 96222 173216 96228
rect 169668 96212 169720 96218
rect 169668 96154 169720 96160
rect 165528 95872 165580 95878
rect 165528 95814 165580 95820
rect 162768 95192 162820 95198
rect 162768 95134 162820 95140
rect 162780 6914 162808 95134
rect 164148 92268 164200 92274
rect 164148 92210 164200 92216
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 153108 3596 153160 3602
rect 153108 3538 153160 3544
rect 154212 3596 154264 3602
rect 154212 3538 154264 3544
rect 155224 3596 155276 3602
rect 155224 3538 155276 3544
rect 155408 3596 155460 3602
rect 155408 3538 155460 3544
rect 155868 3596 155920 3602
rect 155868 3538 155920 3544
rect 156604 3596 156656 3602
rect 156604 3538 156656 3544
rect 157248 3596 157300 3602
rect 157248 3538 157300 3544
rect 157800 3596 157852 3602
rect 157800 3538 157852 3544
rect 158628 3596 158680 3602
rect 158628 3538 158680 3544
rect 158904 3596 158956 3602
rect 158904 3538 158956 3544
rect 160008 3596 160060 3602
rect 160008 3538 160060 3544
rect 160100 3596 160152 3602
rect 160100 3538 160152 3544
rect 161204 3596 161256 3602
rect 161204 3538 161256 3544
rect 154224 480 154252 3538
rect 155420 480 155448 3538
rect 156616 480 156644 3538
rect 157812 480 157840 3538
rect 158916 480 158944 3538
rect 160112 480 160140 3538
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 164160 3602 164188 92210
rect 165540 3602 165568 95814
rect 166908 94444 166960 94450
rect 166908 94386 166960 94392
rect 166920 3602 166948 94386
rect 169024 92336 169076 92342
rect 169024 92278 169076 92284
rect 169036 3602 169064 92278
rect 163688 3596 163740 3602
rect 163688 3538 163740 3544
rect 164148 3596 164200 3602
rect 164148 3538 164200 3544
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 165528 3596 165580 3602
rect 165528 3538 165580 3544
rect 166080 3596 166132 3602
rect 166080 3538 166132 3544
rect 166908 3596 166960 3602
rect 166908 3538 166960 3544
rect 167184 3596 167236 3602
rect 167184 3538 167236 3544
rect 169024 3596 169076 3602
rect 169024 3538 169076 3544
rect 163700 480 163728 3538
rect 164896 480 164924 3538
rect 166092 480 166120 3538
rect 167196 480 167224 3538
rect 169576 3324 169628 3330
rect 169576 3266 169628 3272
rect 168380 3256 168432 3262
rect 168380 3198 168432 3204
rect 168392 480 168420 3198
rect 169588 480 169616 3266
rect 169680 3262 169708 96154
rect 170404 93084 170456 93090
rect 170404 93026 170456 93032
rect 170416 3330 170444 93026
rect 170772 13116 170824 13122
rect 170772 13058 170824 13064
rect 170404 3324 170456 3330
rect 170404 3266 170456 3272
rect 169668 3256 169720 3262
rect 169668 3198 169720 3204
rect 170784 480 170812 13058
rect 173176 3602 173204 96222
rect 174544 94308 174596 94314
rect 174544 94250 174596 94256
rect 171968 3596 172020 3602
rect 171968 3538 172020 3544
rect 173164 3596 173216 3602
rect 173164 3538 173216 3544
rect 174268 3596 174320 3602
rect 174268 3538 174320 3544
rect 171980 480 172008 3538
rect 173164 3256 173216 3262
rect 173164 3198 173216 3204
rect 173176 480 173204 3198
rect 174280 480 174308 3538
rect 174556 3262 174584 94250
rect 175188 92404 175240 92410
rect 175188 92346 175240 92352
rect 175200 3602 175228 92346
rect 176580 3602 176608 96290
rect 177948 94240 178000 94246
rect 177948 94182 178000 94188
rect 177856 92472 177908 92478
rect 177856 92414 177908 92420
rect 175188 3596 175240 3602
rect 175188 3538 175240 3544
rect 175464 3596 175516 3602
rect 175464 3538 175516 3544
rect 176568 3596 176620 3602
rect 176568 3538 176620 3544
rect 176660 3596 176712 3602
rect 176660 3538 176712 3544
rect 174544 3256 174596 3262
rect 174544 3198 174596 3204
rect 175476 480 175504 3538
rect 176672 480 176700 3538
rect 177868 480 177896 92414
rect 177960 3602 177988 94182
rect 179340 6914 179368 96358
rect 180708 93016 180760 93022
rect 180708 92958 180760 92964
rect 179064 6886 179368 6914
rect 177948 3596 178000 3602
rect 177948 3538 178000 3544
rect 179064 480 179092 6886
rect 180720 3602 180748 92958
rect 182088 91724 182140 91730
rect 182088 91666 182140 91672
rect 182100 3602 182128 91666
rect 183480 3602 183508 96426
rect 184848 94172 184900 94178
rect 184848 94114 184900 94120
rect 184860 3602 184888 94114
rect 186976 3602 187004 96562
rect 191104 95804 191156 95810
rect 191104 95746 191156 95752
rect 188344 92948 188396 92954
rect 188344 92890 188396 92896
rect 187056 91656 187108 91662
rect 187056 91598 187108 91604
rect 180248 3596 180300 3602
rect 180248 3538 180300 3544
rect 180708 3596 180760 3602
rect 180708 3538 180760 3544
rect 181444 3596 181496 3602
rect 181444 3538 181496 3544
rect 182088 3596 182140 3602
rect 182088 3538 182140 3544
rect 182548 3596 182600 3602
rect 182548 3538 182600 3544
rect 183468 3596 183520 3602
rect 183468 3538 183520 3544
rect 183744 3596 183796 3602
rect 183744 3538 183796 3544
rect 184848 3596 184900 3602
rect 184848 3538 184900 3544
rect 186136 3596 186188 3602
rect 186136 3538 186188 3544
rect 186964 3596 187016 3602
rect 186964 3538 187016 3544
rect 180260 480 180288 3538
rect 181456 480 181484 3538
rect 182560 480 182588 3538
rect 183756 480 183784 3538
rect 184940 3052 184992 3058
rect 184940 2994 184992 3000
rect 184952 480 184980 2994
rect 186148 480 186176 3538
rect 187068 3058 187096 91598
rect 188356 3602 188384 92890
rect 188988 18624 189040 18630
rect 188988 18566 189040 18572
rect 189000 3602 189028 18566
rect 190828 6588 190880 6594
rect 190828 6530 190880 6536
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 188344 3596 188396 3602
rect 188344 3538 188396 3544
rect 188528 3596 188580 3602
rect 188528 3538 188580 3544
rect 188988 3596 189040 3602
rect 188988 3538 189040 3544
rect 189724 3596 189776 3602
rect 189724 3538 189776 3544
rect 187056 3052 187108 3058
rect 187056 2994 187108 3000
rect 187344 480 187372 3538
rect 188540 480 188568 3538
rect 189736 480 189764 3538
rect 190840 480 190868 6530
rect 191116 3602 191144 95746
rect 192496 7682 192524 97038
rect 195244 96960 195296 96966
rect 195244 96902 195296 96908
rect 194508 95600 194560 95606
rect 194508 95542 194560 95548
rect 192484 7676 192536 7682
rect 192484 7618 192536 7624
rect 192576 7676 192628 7682
rect 192576 7618 192628 7624
rect 192588 3602 192616 7618
rect 194416 6656 194468 6662
rect 194416 6598 194468 6604
rect 191104 3596 191156 3602
rect 191104 3538 191156 3544
rect 192024 3596 192076 3602
rect 192024 3538 192076 3544
rect 192576 3596 192628 3602
rect 192576 3538 192628 3544
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 192036 480 192064 3538
rect 193232 480 193260 3538
rect 194428 480 194456 6598
rect 194520 3602 194548 95542
rect 195256 6254 195284 96902
rect 195348 86290 195376 97815
rect 196624 97164 196676 97170
rect 196624 97106 196676 97112
rect 195336 86284 195388 86290
rect 195336 86226 195388 86232
rect 196636 84862 196664 97106
rect 198004 97028 198056 97034
rect 198004 96970 198056 96976
rect 197268 95736 197320 95742
rect 197268 95678 197320 95684
rect 196624 84856 196676 84862
rect 196624 84798 196676 84804
rect 195612 8016 195664 8022
rect 195612 7958 195664 7964
rect 195244 6248 195296 6254
rect 195244 6190 195296 6196
rect 194508 3596 194560 3602
rect 194508 3538 194560 3544
rect 195624 480 195652 7958
rect 197280 3602 197308 95678
rect 198016 47598 198044 96970
rect 199384 96892 199436 96898
rect 199384 96834 199436 96840
rect 198648 94104 198700 94110
rect 198648 94046 198700 94052
rect 198004 47592 198056 47598
rect 198004 47534 198056 47540
rect 198660 3602 198688 94046
rect 199396 86426 199424 96834
rect 200028 95668 200080 95674
rect 200028 95610 200080 95616
rect 199384 86420 199436 86426
rect 199384 86362 199436 86368
rect 199108 8084 199160 8090
rect 199108 8026 199160 8032
rect 196808 3596 196860 3602
rect 196808 3538 196860 3544
rect 197268 3596 197320 3602
rect 197268 3538 197320 3544
rect 197912 3596 197964 3602
rect 197912 3538 197964 3544
rect 198648 3596 198700 3602
rect 198648 3538 198700 3544
rect 196820 480 196848 3538
rect 197924 480 197952 3538
rect 199120 480 199148 8026
rect 200040 4026 200068 95610
rect 200132 4826 200160 100028
rect 200212 97504 200264 97510
rect 200212 97446 200264 97452
rect 200120 4820 200172 4826
rect 200120 4762 200172 4768
rect 200224 4162 200252 97446
rect 200316 4894 200344 100028
rect 200408 100014 200514 100042
rect 200592 100014 200698 100042
rect 200408 4962 200436 100014
rect 200592 6186 200620 100014
rect 200868 97889 200896 100028
rect 200960 100014 201066 100042
rect 201144 100014 201250 100042
rect 200854 97880 200910 97889
rect 200854 97815 200910 97824
rect 200960 97510 200988 100014
rect 200948 97504 201000 97510
rect 200948 97446 201000 97452
rect 201144 84194 201172 100014
rect 201512 93158 201540 100028
rect 201710 100014 201816 100042
rect 201592 98320 201644 98326
rect 201592 98262 201644 98268
rect 201500 93152 201552 93158
rect 201500 93094 201552 93100
rect 201604 86358 201632 98262
rect 201788 89010 201816 100014
rect 201880 98326 201908 100028
rect 201868 98320 201920 98326
rect 201868 98262 201920 98268
rect 201868 96960 201920 96966
rect 201868 96902 201920 96908
rect 201960 96960 202012 96966
rect 201960 96902 202012 96908
rect 201880 96762 201908 96902
rect 201868 96756 201920 96762
rect 201868 96698 201920 96704
rect 201776 89004 201828 89010
rect 201776 88946 201828 88952
rect 201592 86352 201644 86358
rect 201592 86294 201644 86300
rect 200960 84166 201172 84194
rect 200580 6180 200632 6186
rect 200580 6122 200632 6128
rect 200396 4956 200448 4962
rect 200396 4898 200448 4904
rect 200304 4888 200356 4894
rect 200304 4830 200356 4836
rect 200224 4134 200436 4162
rect 200040 3998 200344 4026
rect 200316 480 200344 3998
rect 200408 3466 200436 4134
rect 200960 3534 200988 84166
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 200948 3528 201000 3534
rect 200948 3470 201000 3476
rect 200396 3460 200448 3466
rect 200396 3402 200448 3408
rect 201512 480 201540 3538
rect 201972 3126 202000 96902
rect 202064 94489 202092 100028
rect 202248 98802 202276 100028
rect 202340 100014 202446 100042
rect 202524 100014 202722 100042
rect 202236 98796 202288 98802
rect 202236 98738 202288 98744
rect 202050 94480 202106 94489
rect 202050 94415 202106 94424
rect 202340 87650 202368 100014
rect 202524 96966 202552 100014
rect 202696 97096 202748 97102
rect 202696 97038 202748 97044
rect 202788 97096 202840 97102
rect 202788 97038 202840 97044
rect 202512 96960 202564 96966
rect 202512 96902 202564 96908
rect 202708 96694 202736 97038
rect 202800 96898 202828 97038
rect 202788 96892 202840 96898
rect 202788 96834 202840 96840
rect 202696 96688 202748 96694
rect 202696 96630 202748 96636
rect 202892 95946 202920 100028
rect 203076 98666 203104 100028
rect 203168 100014 203274 100042
rect 203064 98660 203116 98666
rect 203064 98602 203116 98608
rect 202880 95940 202932 95946
rect 202880 95882 202932 95888
rect 202972 95940 203024 95946
rect 202972 95882 203024 95888
rect 202984 91798 203012 95882
rect 202972 91792 203024 91798
rect 202972 91734 203024 91740
rect 203168 89078 203196 100014
rect 203340 97504 203392 97510
rect 203340 97446 203392 97452
rect 203352 97306 203380 97446
rect 203340 97300 203392 97306
rect 203340 97242 203392 97248
rect 203444 97209 203472 100028
rect 203430 97200 203486 97209
rect 203430 97135 203486 97144
rect 203524 96892 203576 96898
rect 203524 96834 203576 96840
rect 203156 89072 203208 89078
rect 203156 89014 203208 89020
rect 203536 87718 203564 96834
rect 203628 94518 203656 100028
rect 203720 100014 203918 100042
rect 203720 95946 203748 100014
rect 204088 96830 204116 100028
rect 204076 96824 204128 96830
rect 204076 96766 204128 96772
rect 203708 95940 203760 95946
rect 203708 95882 203760 95888
rect 203616 94512 203668 94518
rect 203616 94454 203668 94460
rect 203524 87712 203576 87718
rect 203524 87654 203576 87660
rect 202328 87644 202380 87650
rect 202328 87586 202380 87592
rect 202696 8152 202748 8158
rect 202696 8094 202748 8100
rect 201960 3120 202012 3126
rect 201960 3062 202012 3068
rect 202708 480 202736 8094
rect 204272 3670 204300 100028
rect 204364 100014 204470 100042
rect 204364 7614 204392 100014
rect 204640 98734 204668 100028
rect 204732 100014 204838 100042
rect 205008 100014 205114 100042
rect 204628 98728 204680 98734
rect 204628 98670 204680 98676
rect 204732 89146 204760 100014
rect 204720 89140 204772 89146
rect 204720 89082 204772 89088
rect 205008 8974 205036 100014
rect 205284 94586 205312 100028
rect 205468 97102 205496 100028
rect 205456 97096 205508 97102
rect 205456 97038 205508 97044
rect 205272 94580 205324 94586
rect 205272 94522 205324 94528
rect 205652 9042 205680 100028
rect 205836 98870 205864 100028
rect 205824 98864 205876 98870
rect 205824 98806 205876 98812
rect 205732 97572 205784 97578
rect 205732 97514 205784 97520
rect 205744 97102 205772 97514
rect 206020 97374 206048 100028
rect 206008 97368 206060 97374
rect 206008 97310 206060 97316
rect 205732 97096 205784 97102
rect 205732 97038 205784 97044
rect 206296 94654 206324 100028
rect 206480 96762 206508 100028
rect 206664 97510 206692 100028
rect 206756 100014 206862 100042
rect 206652 97504 206704 97510
rect 206652 97446 206704 97452
rect 206468 96756 206520 96762
rect 206468 96698 206520 96704
rect 206284 94648 206336 94654
rect 206284 94590 206336 94596
rect 206756 90370 206784 100014
rect 207032 98938 207060 100028
rect 207020 98932 207072 98938
rect 207020 98874 207072 98880
rect 206928 97300 206980 97306
rect 206928 97242 206980 97248
rect 206940 96558 206968 97242
rect 207216 96898 207244 100028
rect 207204 96892 207256 96898
rect 207204 96834 207256 96840
rect 206928 96552 206980 96558
rect 206928 96494 206980 96500
rect 207492 91866 207520 100028
rect 207676 99006 207704 100028
rect 207860 99210 207888 100028
rect 207952 100014 208058 100042
rect 208136 100014 208242 100042
rect 207848 99204 207900 99210
rect 207848 99146 207900 99152
rect 207664 99000 207716 99006
rect 207664 98942 207716 98948
rect 207480 91860 207532 91866
rect 207480 91802 207532 91808
rect 206744 90364 206796 90370
rect 206744 90306 206796 90312
rect 207952 89714 207980 100014
rect 208136 99374 208164 100014
rect 208044 99346 208164 99374
rect 208044 90438 208072 99346
rect 208124 97368 208176 97374
rect 208124 97310 208176 97316
rect 208136 95878 208164 97310
rect 208412 96694 208440 100028
rect 208702 100014 208808 100042
rect 208492 98320 208544 98326
rect 208492 98262 208544 98268
rect 208400 96688 208452 96694
rect 208400 96630 208452 96636
rect 208124 95872 208176 95878
rect 208124 95814 208176 95820
rect 208504 91934 208532 98262
rect 208584 94580 208636 94586
rect 208584 94522 208636 94528
rect 208492 91928 208544 91934
rect 208492 91870 208544 91876
rect 208032 90432 208084 90438
rect 208032 90374 208084 90380
rect 207308 89686 207980 89714
rect 205640 9036 205692 9042
rect 205640 8978 205692 8984
rect 204996 8968 205048 8974
rect 204996 8910 205048 8916
rect 204352 7608 204404 7614
rect 204352 7550 204404 7556
rect 207308 5030 207336 89686
rect 208596 87854 208624 94522
rect 208584 87848 208636 87854
rect 208584 87790 208636 87796
rect 208584 6180 208636 6186
rect 208584 6122 208636 6128
rect 207296 5024 207348 5030
rect 207296 4966 207348 4972
rect 207388 4820 207440 4826
rect 207388 4762 207440 4768
rect 204260 3664 204312 3670
rect 204260 3606 204312 3612
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 203892 3460 203944 3466
rect 203892 3402 203944 3408
rect 203904 480 203932 3402
rect 205088 3324 205140 3330
rect 205088 3266 205140 3272
rect 205100 480 205128 3266
rect 206204 480 206232 3470
rect 207400 480 207428 4762
rect 208596 480 208624 6122
rect 208780 3738 208808 100014
rect 208872 98326 208900 100028
rect 208860 98320 208912 98326
rect 208860 98262 208912 98268
rect 208952 97708 209004 97714
rect 208952 97650 209004 97656
rect 208964 97238 208992 97650
rect 208860 97232 208912 97238
rect 208860 97174 208912 97180
rect 208952 97232 209004 97238
rect 208952 97174 209004 97180
rect 208872 96966 208900 97174
rect 208860 96960 208912 96966
rect 208860 96902 208912 96908
rect 209056 96614 209084 100028
rect 208964 96586 209084 96614
rect 209148 100014 209254 100042
rect 209332 100014 209438 100042
rect 209516 100014 209622 100042
rect 208964 87922 208992 96586
rect 208952 87916 209004 87922
rect 208952 87858 209004 87864
rect 209148 86954 209176 100014
rect 209332 90506 209360 100014
rect 209516 94586 209544 100014
rect 209504 94580 209556 94586
rect 209504 94522 209556 94528
rect 209320 90500 209372 90506
rect 209320 90442 209372 90448
rect 208964 86926 209176 86954
rect 208964 5098 208992 86926
rect 209780 7608 209832 7614
rect 209780 7550 209832 7556
rect 208952 5092 209004 5098
rect 208952 5034 209004 5040
rect 208768 3732 208820 3738
rect 208768 3674 208820 3680
rect 209792 480 209820 7550
rect 209884 5166 209912 100028
rect 209964 94512 210016 94518
rect 209964 94454 210016 94460
rect 209976 6390 210004 94454
rect 210068 93226 210096 100028
rect 210252 99074 210280 100028
rect 210450 100014 210556 100042
rect 210240 99068 210292 99074
rect 210240 99010 210292 99016
rect 210424 96688 210476 96694
rect 210424 96630 210476 96636
rect 210148 94580 210200 94586
rect 210148 94522 210200 94528
rect 210056 93220 210108 93226
rect 210056 93162 210108 93168
rect 209964 6384 210016 6390
rect 209964 6326 210016 6332
rect 209872 5160 209924 5166
rect 209872 5102 209924 5108
rect 210160 3806 210188 94522
rect 210436 3874 210464 96630
rect 210528 89714 210556 100014
rect 210620 94586 210648 100028
rect 210804 94722 210832 100028
rect 210896 100014 211094 100042
rect 211278 100014 211384 100042
rect 210792 94716 210844 94722
rect 210792 94658 210844 94664
rect 210608 94580 210660 94586
rect 210608 94522 210660 94528
rect 210896 94518 210924 100014
rect 210884 94512 210936 94518
rect 210884 94454 210936 94460
rect 211356 90574 211384 100014
rect 211448 97034 211476 100028
rect 211632 99482 211660 100028
rect 211724 100014 211830 100042
rect 211620 99476 211672 99482
rect 211620 99418 211672 99424
rect 211724 98274 211752 100014
rect 211804 99476 211856 99482
rect 211804 99418 211856 99424
rect 211540 98246 211752 98274
rect 211436 97028 211488 97034
rect 211436 96970 211488 96976
rect 211344 90568 211396 90574
rect 211344 90510 211396 90516
rect 210528 89686 210740 89714
rect 210712 6322 210740 89686
rect 211540 89214 211568 98246
rect 211816 96614 211844 99418
rect 212000 99278 212028 100028
rect 212092 100014 212290 100042
rect 212368 100014 212474 100042
rect 211988 99272 212040 99278
rect 211988 99214 212040 99220
rect 211632 96586 211844 96614
rect 211632 96014 211660 96586
rect 211620 96008 211672 96014
rect 211620 95950 211672 95956
rect 212092 93294 212120 100014
rect 212080 93288 212132 93294
rect 212080 93230 212132 93236
rect 212368 89714 212396 100014
rect 212540 97504 212592 97510
rect 212540 97446 212592 97452
rect 212552 95062 212580 97446
rect 212644 96966 212672 100028
rect 212632 96960 212684 96966
rect 212632 96902 212684 96908
rect 212540 95056 212592 95062
rect 212540 94998 212592 95004
rect 212828 92002 212856 100028
rect 212908 94580 212960 94586
rect 212908 94522 212960 94528
rect 212816 91996 212868 92002
rect 212816 91938 212868 91944
rect 211724 89686 212396 89714
rect 211724 89350 211752 89686
rect 211712 89344 211764 89350
rect 211712 89286 211764 89292
rect 211528 89208 211580 89214
rect 211528 89150 211580 89156
rect 212920 87786 212948 94522
rect 213012 89282 213040 100028
rect 213104 100014 213210 100042
rect 213288 100014 213486 100042
rect 213564 100014 213670 100042
rect 213104 94790 213132 100014
rect 213092 94784 213144 94790
rect 213092 94726 213144 94732
rect 213288 92070 213316 100014
rect 213564 94586 213592 100014
rect 213840 99142 213868 100028
rect 213932 100014 214038 100042
rect 213828 99136 213880 99142
rect 213828 99078 213880 99084
rect 213932 96642 213960 100014
rect 213840 96614 213960 96642
rect 213552 94580 213604 94586
rect 213552 94522 213604 94528
rect 213840 93362 213868 96614
rect 214104 94580 214156 94586
rect 214104 94522 214156 94528
rect 213828 93356 213880 93362
rect 213828 93298 213880 93304
rect 213276 92064 213328 92070
rect 213276 92006 213328 92012
rect 213000 89276 213052 89282
rect 213000 89218 213052 89224
rect 212908 87780 212960 87786
rect 212908 87722 212960 87728
rect 214116 10402 214144 94522
rect 214104 10396 214156 10402
rect 214104 10338 214156 10344
rect 214208 10334 214236 100028
rect 214392 97918 214420 100028
rect 214484 100014 214682 100042
rect 214760 100014 214866 100042
rect 214944 100014 215050 100042
rect 215128 100014 215234 100042
rect 215418 100014 215524 100042
rect 214380 97912 214432 97918
rect 214380 97854 214432 97860
rect 214484 94568 214512 100014
rect 214760 94586 214788 100014
rect 214300 94540 214512 94568
rect 214748 94580 214800 94586
rect 214196 10328 214248 10334
rect 214196 10270 214248 10276
rect 214300 9110 214328 94540
rect 214748 94522 214800 94528
rect 214944 90642 214972 100014
rect 215128 99374 215156 100014
rect 215036 99346 215156 99374
rect 214932 90636 214984 90642
rect 214932 90578 214984 90584
rect 215036 90522 215064 99346
rect 215300 97912 215352 97918
rect 215300 97854 215352 97860
rect 215116 97844 215168 97850
rect 215116 97786 215168 97792
rect 214484 90494 215064 90522
rect 214484 9178 214512 90494
rect 215128 89714 215156 97786
rect 215312 96082 215340 97854
rect 215496 96914 215524 100014
rect 215588 97442 215616 100028
rect 215576 97436 215628 97442
rect 215576 97378 215628 97384
rect 215760 96960 215812 96966
rect 215496 96886 215708 96914
rect 215760 96902 215812 96908
rect 215484 96824 215536 96830
rect 215484 96766 215536 96772
rect 215300 96076 215352 96082
rect 215300 96018 215352 96024
rect 214668 89686 215156 89714
rect 214668 84194 214696 89686
rect 214576 84166 214696 84194
rect 214472 9172 214524 9178
rect 214472 9114 214524 9120
rect 214288 9104 214340 9110
rect 214288 9046 214340 9052
rect 210700 6316 210752 6322
rect 210700 6258 210752 6264
rect 212172 6248 212224 6254
rect 212172 6190 212224 6196
rect 210976 4888 211028 4894
rect 210976 4830 211028 4836
rect 210424 3868 210476 3874
rect 210424 3810 210476 3816
rect 210148 3800 210200 3806
rect 210148 3742 210200 3748
rect 210988 480 211016 4830
rect 212184 480 212212 6190
rect 214472 4956 214524 4962
rect 214472 4898 214524 4904
rect 213368 3664 213420 3670
rect 213368 3606 213420 3612
rect 213380 480 213408 3606
rect 214484 480 214512 4898
rect 214576 4010 214604 84166
rect 215496 10606 215524 96766
rect 215484 10600 215536 10606
rect 215484 10542 215536 10548
rect 215680 10470 215708 96886
rect 215668 10464 215720 10470
rect 215668 10406 215720 10412
rect 215772 9314 215800 96902
rect 215760 9308 215812 9314
rect 215760 9250 215812 9256
rect 215864 9246 215892 100028
rect 216048 10538 216076 100028
rect 216232 96694 216260 100028
rect 216324 100014 216430 100042
rect 216508 100014 216614 100042
rect 216324 96966 216352 100014
rect 216312 96960 216364 96966
rect 216312 96902 216364 96908
rect 216508 96830 216536 100014
rect 216680 97776 216732 97782
rect 216680 97718 216732 97724
rect 216496 96824 216548 96830
rect 216496 96766 216548 96772
rect 216220 96688 216272 96694
rect 216220 96630 216272 96636
rect 216692 94382 216720 97718
rect 216784 97646 216812 100028
rect 216772 97640 216824 97646
rect 216772 97582 216824 97588
rect 216864 96960 216916 96966
rect 216864 96902 216916 96908
rect 216680 94376 216732 94382
rect 216680 94318 216732 94324
rect 216876 89418 216904 96902
rect 217060 92138 217088 100028
rect 217152 100014 217258 100042
rect 217152 96966 217180 100014
rect 217140 96960 217192 96966
rect 217140 96902 217192 96908
rect 217140 96824 217192 96830
rect 217140 96766 217192 96772
rect 217048 92132 217100 92138
rect 217048 92074 217100 92080
rect 216864 89412 216916 89418
rect 216864 89354 216916 89360
rect 217152 15910 217180 96766
rect 217324 90364 217376 90370
rect 217324 90306 217376 90312
rect 217140 15904 217192 15910
rect 217140 15846 217192 15852
rect 216036 10532 216088 10538
rect 216036 10474 216088 10480
rect 215852 9240 215904 9246
rect 215852 9182 215904 9188
rect 215668 6316 215720 6322
rect 215668 6258 215720 6264
rect 214564 4004 214616 4010
rect 214564 3946 214616 3952
rect 215680 480 215708 6258
rect 216864 3732 216916 3738
rect 216864 3674 216916 3680
rect 216876 480 216904 3674
rect 217336 3330 217364 90306
rect 217428 86494 217456 100028
rect 217520 100014 217626 100042
rect 217704 100014 217810 100042
rect 217520 90710 217548 100014
rect 217704 96830 217732 100014
rect 217980 97170 218008 100028
rect 218060 97436 218112 97442
rect 218060 97378 218112 97384
rect 217968 97164 218020 97170
rect 217968 97106 218020 97112
rect 217692 96824 217744 96830
rect 217692 96766 217744 96772
rect 218072 95606 218100 97378
rect 218256 96830 218284 100028
rect 218348 100014 218454 100042
rect 218244 96824 218296 96830
rect 218244 96766 218296 96772
rect 218060 95600 218112 95606
rect 218060 95542 218112 95548
rect 217508 90704 217560 90710
rect 217508 90646 217560 90652
rect 218348 87990 218376 100014
rect 218520 98388 218572 98394
rect 218520 98330 218572 98336
rect 218532 89486 218560 98330
rect 218624 97578 218652 100028
rect 218822 100014 218928 100042
rect 218900 98274 218928 100014
rect 218992 98394 219020 100028
rect 218980 98388 219032 98394
rect 218980 98330 219032 98336
rect 218900 98246 219112 98274
rect 218612 97572 218664 97578
rect 218612 97514 218664 97520
rect 218796 97572 218848 97578
rect 218796 97514 218848 97520
rect 218808 93702 218836 97514
rect 218888 96824 218940 96830
rect 218888 96766 218940 96772
rect 218796 93696 218848 93702
rect 218796 93638 218848 93644
rect 218900 90778 218928 96766
rect 219084 90846 219112 98246
rect 219176 97102 219204 100028
rect 219164 97096 219216 97102
rect 219164 97038 219216 97044
rect 219452 96830 219480 100028
rect 219650 100014 219756 100042
rect 219728 97170 219756 100014
rect 219820 97850 219848 100028
rect 219912 100014 220018 100042
rect 220096 100014 220202 100042
rect 220280 100014 220386 100042
rect 220464 100014 220662 100042
rect 220846 100014 220952 100042
rect 219808 97844 219860 97850
rect 219808 97786 219860 97792
rect 219716 97164 219768 97170
rect 219716 97106 219768 97112
rect 219912 97050 219940 100014
rect 219544 97022 219940 97050
rect 219440 96824 219492 96830
rect 219440 96766 219492 96772
rect 219072 90840 219124 90846
rect 219072 90782 219124 90788
rect 218888 90772 218940 90778
rect 218888 90714 218940 90720
rect 218520 89480 218572 89486
rect 218520 89422 218572 89428
rect 218336 87984 218388 87990
rect 218336 87926 218388 87932
rect 217416 86488 217468 86494
rect 217416 86430 217468 86436
rect 219544 9450 219572 97022
rect 219716 96960 219768 96966
rect 220096 96948 220124 100014
rect 219716 96902 219768 96908
rect 219912 96920 220124 96948
rect 219728 9518 219756 96902
rect 219912 11762 219940 96920
rect 220280 96778 220308 100014
rect 220360 97164 220412 97170
rect 220360 97106 220412 97112
rect 220096 96750 220308 96778
rect 219900 11756 219952 11762
rect 219900 11698 219952 11704
rect 219716 9512 219768 9518
rect 219716 9454 219768 9460
rect 219532 9444 219584 9450
rect 219532 9386 219584 9392
rect 218060 5024 218112 5030
rect 218060 4966 218112 4972
rect 217324 3324 217376 3330
rect 217324 3266 217376 3272
rect 218072 480 218100 4966
rect 220096 3942 220124 96750
rect 220372 84194 220400 97106
rect 220464 96966 220492 100014
rect 220452 96960 220504 96966
rect 220924 96948 220952 100014
rect 221016 97238 221044 100028
rect 221200 97714 221228 100028
rect 221188 97708 221240 97714
rect 221188 97650 221240 97656
rect 221004 97232 221056 97238
rect 221004 97174 221056 97180
rect 220924 96920 221320 96948
rect 220452 96902 220504 96908
rect 220452 96824 220504 96830
rect 220452 96766 220504 96772
rect 221096 96824 221148 96830
rect 221096 96766 221148 96772
rect 220280 84166 220400 84194
rect 220280 10674 220308 84166
rect 220268 10668 220320 10674
rect 220268 10610 220320 10616
rect 220464 9382 220492 96766
rect 220452 9376 220504 9382
rect 220452 9318 220504 9324
rect 220452 8968 220504 8974
rect 220452 8910 220504 8916
rect 220084 3936 220136 3942
rect 220084 3878 220136 3884
rect 219256 3800 219308 3806
rect 219256 3742 219308 3748
rect 219268 480 219296 3742
rect 220464 480 220492 8910
rect 221108 4078 221136 96766
rect 221292 89554 221320 96920
rect 221384 94858 221412 100028
rect 221464 96960 221516 96966
rect 221464 96902 221516 96908
rect 221372 94852 221424 94858
rect 221372 94794 221424 94800
rect 221476 93430 221504 96902
rect 221464 93424 221516 93430
rect 221464 93366 221516 93372
rect 221568 92206 221596 100028
rect 221660 100014 221858 100042
rect 221936 100014 222042 100042
rect 222226 100014 222332 100042
rect 221660 96830 221688 100014
rect 221936 96966 221964 100014
rect 222304 96966 222332 100014
rect 222396 97918 222424 100028
rect 222594 100014 222700 100042
rect 222384 97912 222436 97918
rect 222384 97854 222436 97860
rect 221924 96960 221976 96966
rect 221924 96902 221976 96908
rect 222292 96960 222344 96966
rect 222292 96902 222344 96908
rect 222476 96892 222528 96898
rect 222476 96834 222528 96840
rect 221648 96824 221700 96830
rect 221648 96766 221700 96772
rect 222292 96824 222344 96830
rect 222292 96766 222344 96772
rect 221556 92200 221608 92206
rect 221556 92142 221608 92148
rect 221280 89548 221332 89554
rect 221280 89490 221332 89496
rect 222304 6526 222332 96766
rect 222488 7886 222516 96834
rect 222476 7880 222528 7886
rect 222476 7822 222528 7828
rect 222292 6520 222344 6526
rect 222292 6462 222344 6468
rect 222672 6458 222700 100014
rect 222764 7818 222792 100028
rect 222936 96960 222988 96966
rect 222936 96902 222988 96908
rect 222752 7812 222804 7818
rect 222752 7754 222804 7760
rect 222948 7750 222976 96902
rect 223040 94926 223068 100028
rect 223132 100014 223238 100042
rect 223316 100014 223422 100042
rect 223132 96830 223160 100014
rect 223316 96898 223344 100014
rect 223304 96892 223356 96898
rect 223304 96834 223356 96840
rect 223120 96824 223172 96830
rect 223120 96766 223172 96772
rect 223028 94920 223080 94926
rect 223028 94862 223080 94868
rect 222936 7744 222988 7750
rect 222936 7686 222988 7692
rect 222660 6452 222712 6458
rect 222660 6394 222712 6400
rect 221556 5092 221608 5098
rect 221556 5034 221608 5040
rect 221096 4072 221148 4078
rect 221096 4014 221148 4020
rect 221568 480 221596 5034
rect 223592 4146 223620 100028
rect 223684 100014 223790 100042
rect 223684 93498 223712 100014
rect 223672 93492 223724 93498
rect 223672 93434 223724 93440
rect 223960 7954 223988 100028
rect 224236 97510 224264 100028
rect 224328 100014 224434 100042
rect 224512 100014 224618 100042
rect 224224 97504 224276 97510
rect 224224 97446 224276 97452
rect 224328 96948 224356 100014
rect 224052 96920 224356 96948
rect 224052 93566 224080 96920
rect 224040 93560 224092 93566
rect 224040 93502 224092 93508
rect 224512 90914 224540 100014
rect 224788 94994 224816 100028
rect 224972 97578 225000 100028
rect 225156 97986 225184 100028
rect 225248 100014 225354 100042
rect 225432 100014 225630 100042
rect 225708 100014 225814 100042
rect 225144 97980 225196 97986
rect 225144 97922 225196 97928
rect 224960 97572 225012 97578
rect 224960 97514 225012 97520
rect 224776 94988 224828 94994
rect 224776 94930 224828 94936
rect 224868 94512 224920 94518
rect 224868 94454 224920 94460
rect 224500 90908 224552 90914
rect 224500 90850 224552 90856
rect 223948 7948 224000 7954
rect 223948 7890 224000 7896
rect 223580 4140 223632 4146
rect 223580 4082 223632 4088
rect 223764 4004 223816 4010
rect 223764 3946 223816 3952
rect 223776 3602 223804 3946
rect 223764 3596 223816 3602
rect 223764 3538 223816 3544
rect 224880 3534 224908 94454
rect 225144 3868 225196 3874
rect 225144 3810 225196 3816
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 224868 3528 224920 3534
rect 224868 3470 224920 3476
rect 222752 3256 222804 3262
rect 222752 3198 222804 3204
rect 222764 480 222792 3198
rect 223960 480 223988 3470
rect 225156 480 225184 3810
rect 225248 3398 225276 100014
rect 225432 93634 225460 100014
rect 225420 93628 225472 93634
rect 225420 93570 225472 93576
rect 225708 90982 225736 100014
rect 225984 96150 226012 100028
rect 226076 100014 226182 100042
rect 225972 96144 226024 96150
rect 225972 96086 226024 96092
rect 226076 93770 226104 100014
rect 226352 97782 226380 100028
rect 226340 97776 226392 97782
rect 226340 97718 226392 97724
rect 226536 95130 226564 100028
rect 226524 95124 226576 95130
rect 226524 95066 226576 95072
rect 226812 93838 226840 100028
rect 226904 100014 227010 100042
rect 226800 93832 226852 93838
rect 226800 93774 226852 93780
rect 226064 93764 226116 93770
rect 226064 93706 226116 93712
rect 225696 90976 225748 90982
rect 225696 90918 225748 90924
rect 226904 89714 226932 100014
rect 227180 97306 227208 100028
rect 227168 97300 227220 97306
rect 227168 97242 227220 97248
rect 227364 95198 227392 100028
rect 227456 100014 227562 100042
rect 227746 100014 227852 100042
rect 227352 95192 227404 95198
rect 227352 95134 227404 95140
rect 227456 92274 227484 100014
rect 227720 97708 227772 97714
rect 227720 97650 227772 97656
rect 227628 97300 227680 97306
rect 227628 97242 227680 97248
rect 227444 92268 227496 92274
rect 227444 92210 227496 92216
rect 226628 89686 226932 89714
rect 226628 14482 226656 89686
rect 226616 14476 226668 14482
rect 226616 14418 226668 14424
rect 227640 6914 227668 97242
rect 227732 96354 227760 97650
rect 227824 97374 227852 100014
rect 227812 97368 227864 97374
rect 227812 97310 227864 97316
rect 227720 96348 227772 96354
rect 227720 96290 227772 96296
rect 228008 94450 228036 100028
rect 227996 94444 228048 94450
rect 227996 94386 228048 94392
rect 228192 92342 228220 100028
rect 228376 96218 228404 100028
rect 228468 100014 228574 100042
rect 228652 100014 228758 100042
rect 228364 96212 228416 96218
rect 228364 96154 228416 96160
rect 228468 93090 228496 100014
rect 228652 99374 228680 100014
rect 228560 99346 228680 99374
rect 228456 93084 228508 93090
rect 228456 93026 228508 93032
rect 228180 92336 228232 92342
rect 228180 92278 228232 92284
rect 228560 92154 228588 99346
rect 228928 96286 228956 100028
rect 228916 96280 228968 96286
rect 228916 96222 228968 96228
rect 228640 95260 228692 95266
rect 228640 95202 228692 95208
rect 228100 92126 228588 92154
rect 228100 13122 228128 92126
rect 228652 89714 228680 95202
rect 229204 94314 229232 100028
rect 229192 94308 229244 94314
rect 229192 94250 229244 94256
rect 229388 92410 229416 100028
rect 229572 97714 229600 100028
rect 229664 100014 229770 100042
rect 229560 97708 229612 97714
rect 229560 97650 229612 97656
rect 229664 94246 229692 100014
rect 229744 94716 229796 94722
rect 229744 94658 229796 94664
rect 229652 94240 229704 94246
rect 229652 94182 229704 94188
rect 229376 92404 229428 92410
rect 229376 92346 229428 92352
rect 228376 89686 228680 89714
rect 228088 13116 228140 13122
rect 228088 13058 228140 13064
rect 227548 6886 227668 6914
rect 226340 3936 226392 3942
rect 226340 3878 226392 3884
rect 225236 3392 225288 3398
rect 225236 3334 225288 3340
rect 226352 480 226380 3878
rect 227548 480 227576 6886
rect 228376 4010 228404 89686
rect 228732 4140 228784 4146
rect 228732 4082 228784 4088
rect 228364 4004 228416 4010
rect 228364 3946 228416 3952
rect 228744 480 228772 4082
rect 229756 3262 229784 94658
rect 229836 92608 229888 92614
rect 229836 92550 229888 92556
rect 229848 3738 229876 92550
rect 229940 92478 229968 100028
rect 230124 96422 230152 100028
rect 230216 100014 230414 100042
rect 230598 100014 230704 100042
rect 230112 96416 230164 96422
rect 230112 96358 230164 96364
rect 230216 93022 230244 100014
rect 230204 93016 230256 93022
rect 230204 92958 230256 92964
rect 229928 92472 229980 92478
rect 229928 92414 229980 92420
rect 230388 91792 230440 91798
rect 230388 91734 230440 91740
rect 229928 3868 229980 3874
rect 229928 3810 229980 3816
rect 229836 3732 229888 3738
rect 229836 3674 229888 3680
rect 229940 3482 229968 3810
rect 230400 3534 230428 91734
rect 230676 91730 230704 100014
rect 230768 96490 230796 100028
rect 230860 100014 230966 100042
rect 231044 100014 231150 100042
rect 230756 96484 230808 96490
rect 230756 96426 230808 96432
rect 230860 94602 230888 100014
rect 230768 94574 230888 94602
rect 230768 94178 230796 94574
rect 230848 94444 230900 94450
rect 230848 94386 230900 94392
rect 230756 94172 230808 94178
rect 230756 94114 230808 94120
rect 230664 91724 230716 91730
rect 230664 91666 230716 91672
rect 230860 18630 230888 94386
rect 231044 91662 231072 100014
rect 231320 96626 231348 100028
rect 231412 100014 231610 100042
rect 231688 100014 231794 100042
rect 231308 96620 231360 96626
rect 231308 96562 231360 96568
rect 231124 94376 231176 94382
rect 231124 94318 231176 94324
rect 231032 91656 231084 91662
rect 231032 91598 231084 91604
rect 230848 18624 230900 18630
rect 230848 18566 230900 18572
rect 231136 3806 231164 94318
rect 231412 92954 231440 100014
rect 231584 96824 231636 96830
rect 231584 96766 231636 96772
rect 231400 92948 231452 92954
rect 231400 92890 231452 92896
rect 231216 92540 231268 92546
rect 231216 92482 231268 92488
rect 231124 3800 231176 3806
rect 231124 3742 231176 3748
rect 231228 3670 231256 92482
rect 231596 89714 231624 96766
rect 231688 94450 231716 100014
rect 231860 97164 231912 97170
rect 231860 97106 231912 97112
rect 231872 94518 231900 97106
rect 231964 95810 231992 100028
rect 232056 100026 232162 100042
rect 232044 100020 232162 100026
rect 232096 100014 232162 100020
rect 232240 100014 232346 100042
rect 232044 99962 232096 99968
rect 232240 96614 232268 100014
rect 232320 99952 232372 99958
rect 232320 99894 232372 99900
rect 232056 96586 232268 96614
rect 231952 95804 232004 95810
rect 231952 95746 232004 95752
rect 231860 94512 231912 94518
rect 231860 94454 231912 94460
rect 231676 94444 231728 94450
rect 231676 94386 231728 94392
rect 231320 89686 231624 89714
rect 231320 8974 231348 89686
rect 231308 8968 231360 8974
rect 231308 8910 231360 8916
rect 232056 7682 232084 96586
rect 232228 91044 232280 91050
rect 232228 90986 232280 90992
rect 232044 7676 232096 7682
rect 232044 7618 232096 7624
rect 232240 6662 232268 90986
rect 232332 89714 232360 99894
rect 232516 97442 232544 100028
rect 232608 100014 232806 100042
rect 232884 100014 232990 100042
rect 232504 97436 232556 97442
rect 232504 97378 232556 97384
rect 232608 91050 232636 100014
rect 232596 91044 232648 91050
rect 232596 90986 232648 90992
rect 232332 89686 232452 89714
rect 232228 6656 232280 6662
rect 232228 6598 232280 6604
rect 232424 6594 232452 89686
rect 232884 84194 232912 100014
rect 233160 95742 233188 100028
rect 233252 100014 233358 100042
rect 233542 100014 233648 100042
rect 233726 100014 233924 100042
rect 233148 95736 233200 95742
rect 233148 95678 233200 95684
rect 233148 95396 233200 95402
rect 233148 95338 233200 95344
rect 232700 84166 232912 84194
rect 232700 8022 232728 84166
rect 232688 8016 232740 8022
rect 232688 7958 232740 7964
rect 232412 6588 232464 6594
rect 232412 6530 232464 6536
rect 231216 3664 231268 3670
rect 231216 3606 231268 3612
rect 233160 3534 233188 95338
rect 233252 94110 233280 100014
rect 233620 99374 233648 100014
rect 233620 99346 233832 99374
rect 233608 94580 233660 94586
rect 233608 94522 233660 94528
rect 233240 94104 233292 94110
rect 233240 94046 233292 94052
rect 233424 91724 233476 91730
rect 233424 91666 233476 91672
rect 233436 8158 233464 91666
rect 233424 8152 233476 8158
rect 233424 8094 233476 8100
rect 229848 3454 229968 3482
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 232228 3528 232280 3534
rect 232228 3470 232280 3476
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 229744 3256 229796 3262
rect 229744 3198 229796 3204
rect 229848 480 229876 3454
rect 231044 480 231072 3470
rect 232240 480 232268 3470
rect 233620 3466 233648 94522
rect 233804 8090 233832 99346
rect 233896 95674 233924 100014
rect 233884 95668 233936 95674
rect 233884 95610 233936 95616
rect 233988 95266 234016 100028
rect 234080 100014 234186 100042
rect 234264 100014 234370 100042
rect 234448 100014 234554 100042
rect 233976 95260 234028 95266
rect 233976 95202 234028 95208
rect 234080 91730 234108 100014
rect 234264 94586 234292 100014
rect 234448 99374 234476 100014
rect 234356 99346 234476 99374
rect 234252 94580 234304 94586
rect 234252 94522 234304 94528
rect 234068 91724 234120 91730
rect 234068 91666 234120 91672
rect 234356 90370 234384 99346
rect 234620 97844 234672 97850
rect 234620 97786 234672 97792
rect 234632 97050 234660 97786
rect 234540 97022 234660 97050
rect 234436 95328 234488 95334
rect 234436 95270 234488 95276
rect 234344 90364 234396 90370
rect 234344 90306 234396 90312
rect 233792 8084 233844 8090
rect 233792 8026 233844 8032
rect 234448 3466 234476 95270
rect 233608 3460 233660 3466
rect 233608 3402 233660 3408
rect 234436 3460 234488 3466
rect 234436 3402 234488 3408
rect 234540 3058 234568 97022
rect 234724 96966 234752 100028
rect 234816 100014 234922 100042
rect 235000 100014 235198 100042
rect 235276 100014 235382 100042
rect 234712 96960 234764 96966
rect 234712 96902 234764 96908
rect 234620 96892 234672 96898
rect 234620 96834 234672 96840
rect 234632 92546 234660 96834
rect 234620 92540 234672 92546
rect 234620 92482 234672 92488
rect 234620 5568 234672 5574
rect 234620 5510 234672 5516
rect 233424 3052 233476 3058
rect 233424 2994 233476 3000
rect 234528 3052 234580 3058
rect 234528 2994 234580 3000
rect 233436 480 233464 2994
rect 234632 480 234660 5510
rect 234816 4826 234844 100014
rect 235000 6186 235028 100014
rect 235276 84194 235304 100014
rect 235448 96960 235500 96966
rect 235448 96902 235500 96908
rect 235092 84166 235304 84194
rect 235092 7614 235120 84166
rect 235080 7608 235132 7614
rect 235080 7550 235132 7556
rect 234988 6180 235040 6186
rect 234988 6122 235040 6128
rect 234804 4820 234856 4826
rect 234804 4762 234856 4768
rect 235460 3602 235488 96902
rect 235552 4894 235580 100028
rect 235644 100014 235750 100042
rect 235828 100014 235934 100042
rect 236118 100014 236224 100042
rect 235644 6254 235672 100014
rect 235828 96898 235856 100014
rect 235816 96892 235868 96898
rect 235816 96834 235868 96840
rect 235632 6248 235684 6254
rect 235632 6190 235684 6196
rect 236196 4962 236224 100014
rect 236288 100014 236394 100042
rect 236288 6322 236316 100014
rect 236460 96960 236512 96966
rect 236460 96902 236512 96908
rect 236276 6316 236328 6322
rect 236276 6258 236328 6264
rect 236472 5098 236500 96902
rect 236564 92614 236592 100028
rect 236656 100014 236762 100042
rect 236552 92608 236604 92614
rect 236552 92550 236604 92556
rect 236460 5092 236512 5098
rect 236460 5034 236512 5040
rect 236656 5030 236684 100014
rect 236932 94382 236960 100028
rect 237116 96830 237144 100028
rect 237208 100014 237314 100042
rect 237208 96966 237236 100014
rect 237196 96960 237248 96966
rect 237196 96902 237248 96908
rect 237104 96824 237156 96830
rect 237104 96766 237156 96772
rect 237576 94722 237604 100028
rect 237760 97170 237788 100028
rect 237748 97164 237800 97170
rect 237748 97106 237800 97112
rect 237656 96960 237708 96966
rect 237656 96902 237708 96908
rect 237564 94716 237616 94722
rect 237564 94658 237616 94664
rect 236920 94376 236972 94382
rect 236920 94318 236972 94324
rect 236644 5024 236696 5030
rect 236644 4966 236696 4972
rect 236184 4956 236236 4962
rect 236184 4898 236236 4904
rect 235540 4888 235592 4894
rect 235540 4830 235592 4836
rect 237668 4146 237696 96902
rect 237656 4140 237708 4146
rect 237656 4082 237708 4088
rect 237944 3942 237972 100028
rect 238142 100014 238248 100042
rect 238116 97980 238168 97986
rect 238116 97922 238168 97928
rect 238024 97912 238076 97918
rect 238024 97854 238076 97860
rect 237932 3936 237984 3942
rect 237932 3878 237984 3884
rect 235448 3596 235500 3602
rect 235448 3538 235500 3544
rect 237012 3460 237064 3466
rect 237012 3402 237064 3408
rect 235816 3188 235868 3194
rect 235816 3130 235868 3136
rect 235828 480 235856 3130
rect 237024 480 237052 3402
rect 238036 3194 238064 97854
rect 238128 3874 238156 97922
rect 238220 4078 238248 100014
rect 238312 97306 238340 100028
rect 238404 100014 238510 100042
rect 238300 97300 238352 97306
rect 238300 97242 238352 97248
rect 238404 96966 238432 100014
rect 238772 97986 238800 100028
rect 238970 100014 239076 100042
rect 238760 97980 238812 97986
rect 238760 97922 238812 97928
rect 239048 96966 239076 100014
rect 238392 96960 238444 96966
rect 238392 96902 238444 96908
rect 239036 96960 239088 96966
rect 239036 96902 239088 96908
rect 239140 95402 239168 100028
rect 239324 97850 239352 100028
rect 239416 100014 239522 100042
rect 239312 97844 239364 97850
rect 239312 97786 239364 97792
rect 239416 97050 239444 100014
rect 239692 97918 239720 100028
rect 239680 97912 239732 97918
rect 239680 97854 239732 97860
rect 239232 97022 239444 97050
rect 239128 95396 239180 95402
rect 239128 95338 239180 95344
rect 239232 84194 239260 97022
rect 239404 96960 239456 96966
rect 239404 96902 239456 96908
rect 239416 91798 239444 96902
rect 239968 95334 239996 100028
rect 240166 100014 240272 100042
rect 240048 97164 240100 97170
rect 240048 97106 240100 97112
rect 239956 95328 240008 95334
rect 239956 95270 240008 95276
rect 239404 91792 239456 91798
rect 239404 91734 239456 91740
rect 239048 84166 239260 84194
rect 239048 5574 239076 84166
rect 240060 15910 240088 97106
rect 240244 96898 240272 100014
rect 240336 96966 240364 100028
rect 240428 100014 240534 100042
rect 240324 96960 240376 96966
rect 240324 96902 240376 96908
rect 240232 96892 240284 96898
rect 240232 96834 240284 96840
rect 240428 84194 240456 100014
rect 240704 96830 240732 100028
rect 240902 100014 241100 100042
rect 241178 100014 241284 100042
rect 240784 96960 240836 96966
rect 240784 96902 240836 96908
rect 240692 96824 240744 96830
rect 240692 96766 240744 96772
rect 240152 84166 240456 84194
rect 240048 15904 240100 15910
rect 240048 15846 240100 15852
rect 239036 5568 239088 5574
rect 239036 5510 239088 5516
rect 238208 4072 238260 4078
rect 238208 4014 238260 4020
rect 238116 3868 238168 3874
rect 238116 3810 238168 3816
rect 238116 3664 238168 3670
rect 238116 3606 238168 3612
rect 238024 3188 238076 3194
rect 238024 3130 238076 3136
rect 238128 480 238156 3606
rect 239312 3188 239364 3194
rect 239312 3130 239364 3136
rect 239324 480 239352 3130
rect 240152 490 240180 84166
rect 240796 3194 240824 96902
rect 240968 96892 241020 96898
rect 240968 96834 241020 96840
rect 240980 3670 241008 96834
rect 241072 93854 241100 100014
rect 241256 96948 241284 100014
rect 241348 97102 241376 100028
rect 241336 97096 241388 97102
rect 241336 97038 241388 97044
rect 241532 96966 241560 100028
rect 241716 97034 241744 100028
rect 241704 97028 241756 97034
rect 241704 96970 241756 96976
rect 241520 96960 241572 96966
rect 241256 96920 241468 96948
rect 241336 96824 241388 96830
rect 241336 96766 241388 96772
rect 241072 93826 241284 93854
rect 241256 4214 241284 93826
rect 241244 4208 241296 4214
rect 241244 4150 241296 4156
rect 240968 3664 241020 3670
rect 240968 3606 241020 3612
rect 241348 3482 241376 96766
rect 241440 3602 241468 96920
rect 241520 96902 241572 96908
rect 241900 96830 241928 100028
rect 242084 97782 242112 100028
rect 242072 97776 242124 97782
rect 242072 97718 242124 97724
rect 242164 97096 242216 97102
rect 242164 97038 242216 97044
rect 241888 96824 241940 96830
rect 241888 96766 241940 96772
rect 241428 3596 241480 3602
rect 241428 3538 241480 3544
rect 241348 3454 241744 3482
rect 240784 3188 240836 3194
rect 240784 3130 240836 3136
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 3454
rect 242176 3262 242204 97038
rect 242360 96898 242388 100028
rect 242558 100014 242664 100042
rect 242532 97028 242584 97034
rect 242532 96970 242584 96976
rect 242440 96960 242492 96966
rect 242440 96902 242492 96908
rect 242348 96892 242400 96898
rect 242348 96834 242400 96840
rect 242452 3330 242480 96902
rect 242440 3324 242492 3330
rect 242440 3266 242492 3272
rect 242164 3256 242216 3262
rect 242164 3198 242216 3204
rect 242544 3126 242572 96970
rect 242636 3738 242664 100014
rect 242728 97170 242756 100028
rect 242716 97164 242768 97170
rect 242716 97106 242768 97112
rect 242808 96892 242860 96898
rect 242808 96834 242860 96840
rect 242716 96824 242768 96830
rect 242716 96766 242768 96772
rect 242624 3732 242676 3738
rect 242624 3674 242676 3680
rect 242728 3398 242756 96766
rect 242820 3874 242848 96834
rect 242912 95742 242940 100028
rect 243096 96694 243124 100028
rect 243280 97374 243308 100028
rect 243570 100014 243676 100042
rect 243268 97368 243320 97374
rect 243268 97310 243320 97316
rect 243084 96688 243136 96694
rect 243084 96630 243136 96636
rect 242900 95736 242952 95742
rect 242900 95678 242952 95684
rect 243648 93226 243676 100014
rect 243740 96966 243768 100028
rect 243728 96960 243780 96966
rect 243728 96902 243780 96908
rect 243636 93220 243688 93226
rect 243636 93162 243688 93168
rect 243924 11762 243952 100028
rect 244016 100014 244122 100042
rect 244016 91798 244044 100014
rect 244096 96960 244148 96966
rect 244096 96902 244148 96908
rect 244004 91792 244056 91798
rect 244004 91734 244056 91740
rect 244108 90370 244136 96902
rect 244292 96762 244320 100028
rect 244476 97442 244504 100028
rect 244464 97436 244516 97442
rect 244464 97378 244516 97384
rect 244752 96966 244780 100028
rect 244740 96960 244792 96966
rect 244740 96902 244792 96908
rect 244280 96756 244332 96762
rect 244280 96698 244332 96704
rect 244936 94654 244964 100028
rect 245134 100014 245240 100042
rect 245108 96892 245160 96898
rect 245108 96834 245160 96840
rect 244924 94648 244976 94654
rect 244924 94590 244976 94596
rect 244096 90364 244148 90370
rect 244096 90306 244148 90312
rect 243912 11756 243964 11762
rect 243912 11698 243964 11704
rect 242900 4208 242952 4214
rect 242900 4150 242952 4156
rect 242808 3868 242860 3874
rect 242808 3810 242860 3816
rect 242716 3392 242768 3398
rect 242716 3334 242768 3340
rect 242532 3120 242584 3126
rect 242532 3062 242584 3068
rect 242912 480 242940 4150
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 244108 480 244136 3538
rect 245120 3534 245148 96834
rect 245212 11830 245240 100014
rect 245200 11824 245252 11830
rect 245200 11766 245252 11772
rect 245304 5030 245332 100028
rect 245384 96960 245436 96966
rect 245384 96902 245436 96908
rect 245396 5234 245424 96902
rect 245488 96898 245516 100028
rect 245476 96892 245528 96898
rect 245476 96834 245528 96840
rect 245672 96830 245700 100028
rect 245948 96966 245976 100028
rect 245936 96960 245988 96966
rect 245936 96902 245988 96908
rect 246132 96898 246160 100028
rect 246316 97306 246344 100028
rect 246304 97300 246356 97306
rect 246304 97242 246356 97248
rect 246120 96892 246172 96898
rect 246120 96834 246172 96840
rect 245660 96824 245712 96830
rect 245660 96766 245712 96772
rect 245476 96756 245528 96762
rect 245476 96698 245528 96704
rect 245384 5228 245436 5234
rect 245384 5170 245436 5176
rect 245292 5024 245344 5030
rect 245292 4966 245344 4972
rect 245488 3602 245516 96698
rect 246304 96688 246356 96694
rect 246304 96630 246356 96636
rect 246316 3670 246344 96630
rect 246500 4962 246528 100028
rect 246684 97102 246712 100028
rect 246776 100014 246882 100042
rect 246672 97096 246724 97102
rect 246672 97038 246724 97044
rect 246580 96960 246632 96966
rect 246776 96948 246804 100014
rect 246856 97096 246908 97102
rect 246856 97038 246908 97044
rect 246580 96902 246632 96908
rect 246684 96920 246804 96948
rect 246488 4956 246540 4962
rect 246488 4898 246540 4904
rect 246304 3664 246356 3670
rect 246304 3606 246356 3612
rect 245476 3596 245528 3602
rect 245476 3538 245528 3544
rect 245108 3528 245160 3534
rect 245108 3470 245160 3476
rect 246592 3466 246620 96902
rect 246684 83502 246712 96920
rect 246764 96824 246816 96830
rect 246764 96766 246816 96772
rect 246672 83496 246724 83502
rect 246672 83438 246724 83444
rect 246776 13122 246804 96766
rect 246868 93158 246896 97038
rect 247144 96966 247172 100028
rect 247328 97714 247356 100028
rect 247316 97708 247368 97714
rect 247316 97650 247368 97656
rect 247512 97578 247540 100028
rect 247500 97572 247552 97578
rect 247500 97514 247552 97520
rect 247132 96960 247184 96966
rect 247132 96902 247184 96908
rect 246948 96892 247000 96898
rect 246948 96834 247000 96840
rect 246856 93152 246908 93158
rect 246856 93094 246908 93100
rect 246960 91866 246988 96834
rect 247696 95946 247724 100028
rect 247894 100014 248000 100042
rect 247684 95940 247736 95946
rect 247684 95882 247736 95888
rect 247972 93854 248000 100014
rect 248064 94586 248092 100028
rect 248156 100014 248354 100042
rect 248052 94580 248104 94586
rect 248052 94522 248104 94528
rect 247972 93826 248092 93854
rect 246948 91860 247000 91866
rect 246948 91802 247000 91808
rect 248064 80714 248092 93826
rect 248156 89010 248184 100014
rect 248420 97436 248472 97442
rect 248420 97378 248472 97384
rect 248432 97238 248460 97378
rect 248420 97232 248472 97238
rect 248420 97174 248472 97180
rect 248524 96966 248552 100028
rect 248236 96960 248288 96966
rect 248236 96902 248288 96908
rect 248512 96960 248564 96966
rect 248512 96902 248564 96908
rect 248144 89004 248196 89010
rect 248144 88946 248196 88952
rect 248248 82142 248276 96902
rect 248708 96898 248736 100028
rect 248906 100014 249012 100042
rect 249090 100014 249196 100042
rect 249274 100014 249472 100042
rect 249550 100014 249656 100042
rect 248696 96892 248748 96898
rect 248696 96834 248748 96840
rect 248984 93854 249012 100014
rect 249168 96914 249196 100014
rect 249340 96960 249392 96966
rect 249168 96886 249288 96914
rect 249340 96902 249392 96908
rect 248984 93826 249196 93854
rect 248236 82136 248288 82142
rect 248236 82078 248288 82084
rect 248052 80708 248104 80714
rect 248052 80650 248104 80656
rect 246764 13116 246816 13122
rect 246764 13058 246816 13064
rect 249168 5166 249196 93826
rect 249260 6186 249288 96886
rect 249352 6730 249380 96902
rect 249340 6724 249392 6730
rect 249340 6666 249392 6672
rect 249248 6180 249300 6186
rect 249248 6122 249300 6128
rect 249156 5160 249208 5166
rect 249156 5102 249208 5108
rect 249444 4826 249472 100014
rect 249524 96892 249576 96898
rect 249524 96834 249576 96840
rect 249536 4894 249564 96834
rect 249628 5098 249656 100014
rect 249720 94518 249748 100028
rect 249904 95606 249932 100028
rect 250088 97034 250116 100028
rect 250076 97028 250128 97034
rect 250076 96970 250128 96976
rect 250272 96898 250300 100028
rect 250456 97646 250484 100028
rect 250444 97640 250496 97646
rect 250444 97582 250496 97588
rect 250640 96966 250668 100028
rect 250720 97028 250772 97034
rect 250720 96970 250772 96976
rect 250628 96960 250680 96966
rect 250628 96902 250680 96908
rect 250260 96892 250312 96898
rect 250260 96834 250312 96840
rect 250444 95736 250496 95742
rect 250444 95678 250496 95684
rect 249892 95600 249944 95606
rect 249892 95542 249944 95548
rect 249708 94512 249760 94518
rect 249708 94454 249760 94460
rect 249984 7608 250036 7614
rect 249984 7550 250036 7556
rect 249616 5092 249668 5098
rect 249616 5034 249668 5040
rect 249524 4888 249576 4894
rect 249524 4830 249576 4836
rect 249432 4820 249484 4826
rect 249432 4762 249484 4768
rect 246580 3460 246632 3466
rect 246580 3402 246632 3408
rect 246396 3324 246448 3330
rect 246396 3266 246448 3272
rect 248788 3324 248840 3330
rect 248788 3266 248840 3272
rect 245200 3256 245252 3262
rect 245200 3198 245252 3204
rect 245212 480 245240 3198
rect 246408 480 246436 3266
rect 247592 3120 247644 3126
rect 247592 3062 247644 3068
rect 247604 480 247632 3062
rect 248800 480 248828 3266
rect 249996 480 250024 7550
rect 250456 3262 250484 95678
rect 250732 6254 250760 96970
rect 250812 96892 250864 96898
rect 250812 96834 250864 96840
rect 250824 16114 250852 96834
rect 250812 16108 250864 16114
rect 250812 16050 250864 16056
rect 250916 16046 250944 100028
rect 250996 96960 251048 96966
rect 250996 96902 251048 96908
rect 250904 16040 250956 16046
rect 250904 15982 250956 15988
rect 251008 10946 251036 96902
rect 251100 95742 251128 100028
rect 251284 97034 251312 100028
rect 251272 97028 251324 97034
rect 251272 96970 251324 96976
rect 251468 96966 251496 100028
rect 251652 97850 251680 100028
rect 251640 97844 251692 97850
rect 251640 97786 251692 97792
rect 251456 96960 251508 96966
rect 251456 96902 251508 96908
rect 251836 96898 251864 100028
rect 252008 96960 252060 96966
rect 252008 96902 252060 96908
rect 251824 96892 251876 96898
rect 251824 96834 251876 96840
rect 251088 95736 251140 95742
rect 251088 95678 251140 95684
rect 250996 10940 251048 10946
rect 250996 10882 251048 10888
rect 250720 6248 250772 6254
rect 250720 6190 250772 6196
rect 251180 3868 251232 3874
rect 251180 3810 251232 3816
rect 250444 3256 250496 3262
rect 250444 3198 250496 3204
rect 251192 480 251220 3810
rect 252020 3806 252048 96902
rect 252112 15978 252140 100028
rect 252296 97034 252324 100028
rect 252388 100014 252494 100042
rect 252192 97028 252244 97034
rect 252192 96970 252244 96976
rect 252284 97028 252336 97034
rect 252284 96970 252336 96976
rect 252100 15972 252152 15978
rect 252100 15914 252152 15920
rect 252204 10878 252232 96970
rect 252284 96892 252336 96898
rect 252284 96834 252336 96840
rect 252192 10872 252244 10878
rect 252192 10814 252244 10820
rect 252296 10810 252324 96834
rect 252284 10804 252336 10810
rect 252284 10746 252336 10752
rect 252388 10742 252416 100014
rect 252468 97028 252520 97034
rect 252468 96970 252520 96976
rect 252480 95810 252508 96970
rect 252664 96966 252692 100028
rect 252652 96960 252704 96966
rect 252652 96902 252704 96908
rect 252468 95804 252520 95810
rect 252468 95746 252520 95752
rect 252848 94246 252876 100028
rect 253032 95878 253060 100028
rect 253322 100014 253428 100042
rect 253296 97776 253348 97782
rect 253296 97718 253348 97724
rect 253204 97708 253256 97714
rect 253204 97650 253256 97656
rect 253020 95872 253072 95878
rect 253020 95814 253072 95820
rect 252836 94240 252888 94246
rect 252836 94182 252888 94188
rect 252376 10736 252428 10742
rect 252376 10678 252428 10684
rect 253216 8974 253244 97650
rect 253308 97374 253336 97718
rect 253296 97368 253348 97374
rect 253296 97310 253348 97316
rect 253400 96914 253428 100014
rect 253492 97102 253520 100028
rect 253584 100014 253690 100042
rect 253480 97096 253532 97102
rect 253480 97038 253532 97044
rect 253400 96886 253520 96914
rect 253388 96824 253440 96830
rect 253388 96766 253440 96772
rect 253400 85474 253428 96766
rect 253388 85468 253440 85474
rect 253388 85410 253440 85416
rect 253492 72486 253520 96886
rect 253584 90098 253612 100014
rect 253756 97096 253808 97102
rect 253756 97038 253808 97044
rect 253664 96960 253716 96966
rect 253664 96902 253716 96908
rect 253572 90092 253624 90098
rect 253572 90034 253624 90040
rect 253676 88806 253704 96902
rect 253768 94314 253796 97038
rect 253860 96830 253888 100028
rect 254044 97714 254072 100028
rect 254032 97708 254084 97714
rect 254032 97650 254084 97656
rect 254228 96966 254256 100028
rect 254518 100014 254624 100042
rect 254216 96960 254268 96966
rect 254216 96902 254268 96908
rect 254596 96914 254624 100014
rect 254688 97034 254716 100028
rect 254886 100014 254992 100042
rect 254676 97028 254728 97034
rect 254676 96970 254728 96976
rect 254596 96886 254900 96914
rect 253848 96824 253900 96830
rect 253848 96766 253900 96772
rect 254768 96824 254820 96830
rect 254768 96766 254820 96772
rect 253756 94308 253808 94314
rect 253756 94250 253808 94256
rect 253664 88800 253716 88806
rect 253664 88742 253716 88748
rect 253480 72480 253532 72486
rect 253480 72422 253532 72428
rect 253480 15904 253532 15910
rect 253480 15846 253532 15852
rect 253204 8968 253256 8974
rect 253204 8910 253256 8916
rect 252008 3800 252060 3806
rect 252008 3742 252060 3748
rect 252376 3732 252428 3738
rect 252376 3674 252428 3680
rect 252388 480 252416 3674
rect 253492 480 253520 15846
rect 254780 6594 254808 96766
rect 254872 15910 254900 96886
rect 254860 15904 254912 15910
rect 254860 15846 254912 15852
rect 254964 10606 254992 100014
rect 255056 97102 255084 100028
rect 255044 97096 255096 97102
rect 255044 97038 255096 97044
rect 255136 97028 255188 97034
rect 255136 96970 255188 96976
rect 255044 96960 255096 96966
rect 255044 96902 255096 96908
rect 255056 10674 255084 96902
rect 255044 10668 255096 10674
rect 255044 10610 255096 10616
rect 254952 10600 255004 10606
rect 254952 10542 255004 10548
rect 255148 6662 255176 96970
rect 255240 96830 255268 100028
rect 255424 96830 255452 100028
rect 255700 96966 255728 100028
rect 255688 96960 255740 96966
rect 255688 96902 255740 96908
rect 255228 96824 255280 96830
rect 255228 96766 255280 96772
rect 255412 96824 255464 96830
rect 255412 96766 255464 96772
rect 255884 94382 255912 100028
rect 256068 97034 256096 100028
rect 256056 97028 256108 97034
rect 256056 96970 256108 96976
rect 256148 96960 256200 96966
rect 256148 96902 256200 96908
rect 256056 96824 256108 96830
rect 256056 96766 256108 96772
rect 255872 94376 255924 94382
rect 255872 94318 255924 94324
rect 256068 91662 256096 96766
rect 256056 91656 256108 91662
rect 256056 91598 256108 91604
rect 255964 90364 256016 90370
rect 255964 90306 256016 90312
rect 255136 6656 255188 6662
rect 255136 6598 255188 6604
rect 254768 6588 254820 6594
rect 254768 6530 254820 6536
rect 255976 3874 256004 90306
rect 256160 86222 256188 96902
rect 256148 86216 256200 86222
rect 256148 86158 256200 86164
rect 256252 13530 256280 100028
rect 256450 100014 256556 100042
rect 256424 97028 256476 97034
rect 256424 96970 256476 96976
rect 256332 96960 256384 96966
rect 256332 96902 256384 96908
rect 256344 90166 256372 96902
rect 256332 90160 256384 90166
rect 256332 90102 256384 90108
rect 256436 88874 256464 96970
rect 256528 92954 256556 100014
rect 256620 96966 256648 100028
rect 256896 98462 256924 100028
rect 256884 98456 256936 98462
rect 256884 98398 256936 98404
rect 256700 97844 256752 97850
rect 256700 97786 256752 97792
rect 256608 96960 256660 96966
rect 256608 96902 256660 96908
rect 256712 95674 256740 97786
rect 256976 97436 257028 97442
rect 256976 97378 257028 97384
rect 256700 95668 256752 95674
rect 256700 95610 256752 95616
rect 256516 92948 256568 92954
rect 256516 92890 256568 92896
rect 256424 88868 256476 88874
rect 256424 88810 256476 88816
rect 256988 16574 257016 97378
rect 257080 96898 257108 100028
rect 257264 97034 257292 100028
rect 257448 97510 257476 100028
rect 257436 97504 257488 97510
rect 257436 97446 257488 97452
rect 257252 97028 257304 97034
rect 257252 96970 257304 96976
rect 257632 96966 257660 100028
rect 257724 100014 257830 100042
rect 257620 96960 257672 96966
rect 257620 96902 257672 96908
rect 257068 96892 257120 96898
rect 257068 96834 257120 96840
rect 257344 93220 257396 93226
rect 257344 93162 257396 93168
rect 256988 16546 257108 16574
rect 256240 13524 256292 13530
rect 256240 13466 256292 13472
rect 256056 11824 256108 11830
rect 256056 11766 256108 11772
rect 256068 3942 256096 11766
rect 256148 11756 256200 11762
rect 256148 11698 256200 11704
rect 256160 4078 256188 11698
rect 256148 4072 256200 4078
rect 256148 4014 256200 4020
rect 256056 3936 256108 3942
rect 256056 3878 256108 3884
rect 255964 3868 256016 3874
rect 255964 3810 256016 3816
rect 255872 3664 255924 3670
rect 255872 3606 255924 3612
rect 254676 3256 254728 3262
rect 254676 3198 254728 3204
rect 254688 480 254716 3198
rect 255884 480 255912 3606
rect 257080 480 257108 16546
rect 257356 4146 257384 93162
rect 257724 88942 257752 100014
rect 258092 97034 258120 100028
rect 257896 97028 257948 97034
rect 257896 96970 257948 96976
rect 258080 97028 258132 97034
rect 258080 96970 258132 96976
rect 257804 96892 257856 96898
rect 257804 96834 257856 96840
rect 257816 93022 257844 96834
rect 257804 93016 257856 93022
rect 257804 92958 257856 92964
rect 257908 90234 257936 96970
rect 257988 96960 258040 96966
rect 257988 96902 258040 96908
rect 258000 93090 258028 96902
rect 258276 96830 258304 100028
rect 258356 97368 258408 97374
rect 258356 97310 258408 97316
rect 258264 96824 258316 96830
rect 258264 96766 258316 96772
rect 258368 93854 258396 97310
rect 258460 96966 258488 100028
rect 258644 98530 258672 100028
rect 258632 98524 258684 98530
rect 258632 98466 258684 98472
rect 258724 97572 258776 97578
rect 258724 97514 258776 97520
rect 258448 96960 258500 96966
rect 258448 96902 258500 96908
rect 258368 93826 258488 93854
rect 257988 93084 258040 93090
rect 257988 93026 258040 93032
rect 257896 90228 257948 90234
rect 257896 90170 257948 90176
rect 257712 88936 257764 88942
rect 257712 88878 257764 88884
rect 258460 7614 258488 93826
rect 258736 14482 258764 97514
rect 258828 96898 258856 100028
rect 259026 100014 259224 100042
rect 259092 97028 259144 97034
rect 259092 96970 259144 96976
rect 259000 96960 259052 96966
rect 259000 96902 259052 96908
rect 258816 96892 258868 96898
rect 258816 96834 258868 96840
rect 259012 89690 259040 96902
rect 259000 89684 259052 89690
rect 259000 89626 259052 89632
rect 259104 85338 259132 96970
rect 259196 96948 259224 100014
rect 259288 97782 259316 100028
rect 259276 97776 259328 97782
rect 259276 97718 259328 97724
rect 259472 96966 259500 100028
rect 259460 96960 259512 96966
rect 259196 96920 259316 96948
rect 259184 96824 259236 96830
rect 259184 96766 259236 96772
rect 259092 85332 259144 85338
rect 259092 85274 259144 85280
rect 258724 14476 258776 14482
rect 258724 14418 258776 14424
rect 258448 7608 258500 7614
rect 258448 7550 258500 7556
rect 259196 6526 259224 96766
rect 259184 6520 259236 6526
rect 259184 6462 259236 6468
rect 257344 4140 257396 4146
rect 257344 4082 257396 4088
rect 258264 4140 258316 4146
rect 258264 4082 258316 4088
rect 258276 480 258304 4082
rect 259288 4010 259316 96920
rect 259460 96902 259512 96908
rect 259656 96898 259684 100028
rect 259368 96892 259420 96898
rect 259368 96834 259420 96840
rect 259644 96892 259696 96898
rect 259644 96834 259696 96840
rect 259276 4004 259328 4010
rect 259276 3946 259328 3952
rect 259380 3806 259408 96834
rect 259840 94450 259868 100028
rect 260024 96762 260052 100028
rect 260104 97232 260156 97238
rect 260104 97174 260156 97180
rect 260012 96756 260064 96762
rect 260012 96698 260064 96704
rect 259828 94444 259880 94450
rect 259828 94386 259880 94392
rect 260116 8294 260144 97174
rect 260208 96830 260236 100028
rect 260484 97374 260512 100028
rect 260576 100014 260682 100042
rect 260472 97368 260524 97374
rect 260472 97310 260524 97316
rect 260288 96960 260340 96966
rect 260576 96948 260604 100014
rect 260288 96902 260340 96908
rect 260392 96920 260604 96948
rect 260196 96824 260248 96830
rect 260196 96766 260248 96772
rect 260104 8288 260156 8294
rect 260104 8230 260156 8236
rect 260300 6458 260328 96902
rect 260288 6452 260340 6458
rect 260288 6394 260340 6400
rect 260392 6322 260420 96920
rect 260748 96892 260800 96898
rect 260748 96834 260800 96840
rect 260472 96824 260524 96830
rect 260472 96766 260524 96772
rect 260484 87582 260512 96766
rect 260564 96756 260616 96762
rect 260564 96698 260616 96704
rect 260472 87576 260524 87582
rect 260472 87518 260524 87524
rect 260576 6390 260604 96698
rect 260760 91730 260788 96834
rect 260852 96694 260880 100028
rect 261036 97170 261064 100028
rect 261024 97164 261076 97170
rect 261024 97106 261076 97112
rect 261220 96966 261248 100028
rect 261208 96960 261260 96966
rect 261208 96902 261260 96908
rect 261404 96762 261432 100028
rect 261680 96898 261708 100028
rect 261878 100014 261984 100042
rect 261760 97028 261812 97034
rect 261760 96970 261812 96976
rect 261668 96892 261720 96898
rect 261668 96834 261720 96840
rect 261392 96756 261444 96762
rect 261392 96698 261444 96704
rect 260840 96688 260892 96694
rect 260840 96630 260892 96636
rect 261484 93152 261536 93158
rect 261484 93094 261536 93100
rect 260748 91724 260800 91730
rect 260748 91666 260800 91672
rect 260564 6384 260616 6390
rect 260564 6326 260616 6332
rect 260380 6316 260432 6322
rect 260380 6258 260432 6264
rect 260656 4072 260708 4078
rect 260656 4014 260708 4020
rect 259460 3868 259512 3874
rect 259460 3810 259512 3816
rect 259368 3800 259420 3806
rect 259368 3742 259420 3748
rect 259472 480 259500 3810
rect 260668 480 260696 4014
rect 261496 3874 261524 93094
rect 261772 86902 261800 96970
rect 261852 96960 261904 96966
rect 261852 96902 261904 96908
rect 261864 93838 261892 96902
rect 261956 96880 261984 100014
rect 262048 97034 262076 100028
rect 262036 97028 262088 97034
rect 262036 96970 262088 96976
rect 261956 96852 262168 96880
rect 262036 96756 262088 96762
rect 262036 96698 262088 96704
rect 261944 96688 261996 96694
rect 261944 96630 261996 96636
rect 261852 93832 261904 93838
rect 261852 93774 261904 93780
rect 261956 88330 261984 96630
rect 261944 88324 261996 88330
rect 261944 88266 261996 88272
rect 262048 88262 262076 96698
rect 262140 93770 262168 96852
rect 262232 96762 262260 100028
rect 262416 96830 262444 100028
rect 262600 97578 262628 100028
rect 262890 100014 262996 100042
rect 262968 97714 262996 100014
rect 263060 98598 263088 100028
rect 263258 100014 263364 100042
rect 263048 98592 263100 98598
rect 263048 98534 263100 98540
rect 262772 97708 262824 97714
rect 262772 97650 262824 97656
rect 262956 97708 263008 97714
rect 262956 97650 263008 97656
rect 262588 97572 262640 97578
rect 262588 97514 262640 97520
rect 262404 96824 262456 96830
rect 262404 96766 262456 96772
rect 262220 96756 262272 96762
rect 262220 96698 262272 96704
rect 262784 94178 262812 97650
rect 262864 97640 262916 97646
rect 262864 97582 262916 97588
rect 262876 95538 262904 97582
rect 263048 97504 263100 97510
rect 263048 97446 263100 97452
rect 262956 96892 263008 96898
rect 262956 96834 263008 96840
rect 262864 95532 262916 95538
rect 262864 95474 262916 95480
rect 262864 94648 262916 94654
rect 262864 94590 262916 94596
rect 262772 94172 262824 94178
rect 262772 94114 262824 94120
rect 262128 93764 262180 93770
rect 262128 93706 262180 93712
rect 262220 91792 262272 91798
rect 262220 91734 262272 91740
rect 262036 88256 262088 88262
rect 262036 88198 262088 88204
rect 261760 86896 261812 86902
rect 261760 86838 261812 86844
rect 261484 3868 261536 3874
rect 261484 3810 261536 3816
rect 262232 3602 262260 91734
rect 262876 3602 262904 94590
rect 262968 83842 262996 96834
rect 263060 85406 263088 97446
rect 263336 96948 263364 100014
rect 263428 97442 263456 100028
rect 263416 97436 263468 97442
rect 263416 97378 263468 97384
rect 263612 97034 263640 100028
rect 263600 97028 263652 97034
rect 263600 96970 263652 96976
rect 263336 96920 263548 96948
rect 263324 96824 263376 96830
rect 263324 96766 263376 96772
rect 263336 93702 263364 96766
rect 263416 96756 263468 96762
rect 263416 96698 263468 96704
rect 263324 93696 263376 93702
rect 263324 93638 263376 93644
rect 263428 90302 263456 96698
rect 263416 90296 263468 90302
rect 263416 90238 263468 90244
rect 263520 88194 263548 96920
rect 263796 96830 263824 100028
rect 264072 96966 264100 100028
rect 264060 96960 264112 96966
rect 264060 96902 264112 96908
rect 264256 96898 264284 100028
rect 264244 96892 264296 96898
rect 264244 96834 264296 96840
rect 263784 96824 263836 96830
rect 263784 96766 263836 96772
rect 264244 91860 264296 91866
rect 264244 91802 264296 91808
rect 263508 88188 263560 88194
rect 263508 88130 263560 88136
rect 263048 85400 263100 85406
rect 263048 85342 263100 85348
rect 262956 83836 263008 83842
rect 262956 83778 263008 83784
rect 264152 8288 264204 8294
rect 264152 8230 264204 8236
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 261760 3596 261812 3602
rect 261760 3538 261812 3544
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 262864 3596 262916 3602
rect 262864 3538 262916 3544
rect 261772 480 261800 3538
rect 262968 480 262996 3606
rect 264164 480 264192 8230
rect 264256 3670 264284 91802
rect 264440 86766 264468 100028
rect 264624 97850 264652 100028
rect 264716 100014 264822 100042
rect 264612 97844 264664 97850
rect 264612 97786 264664 97792
rect 264520 96960 264572 96966
rect 264716 96948 264744 100014
rect 264796 97028 264848 97034
rect 264796 96970 264848 96976
rect 264520 96902 264572 96908
rect 264624 96920 264744 96948
rect 264428 86760 264480 86766
rect 264428 86702 264480 86708
rect 264532 82414 264560 96902
rect 264624 92410 264652 96920
rect 264704 96824 264756 96830
rect 264704 96766 264756 96772
rect 264612 92404 264664 92410
rect 264612 92346 264664 92352
rect 264716 88126 264744 96766
rect 264808 93634 264836 96970
rect 264888 96892 264940 96898
rect 264888 96834 264940 96840
rect 264796 93628 264848 93634
rect 264796 93570 264848 93576
rect 264900 92478 264928 96834
rect 264992 96762 265020 100028
rect 265268 96966 265296 100028
rect 265452 97034 265480 100028
rect 265440 97028 265492 97034
rect 265440 96970 265492 96976
rect 265256 96960 265308 96966
rect 265256 96902 265308 96908
rect 265636 96830 265664 100028
rect 265820 97646 265848 100028
rect 266018 100014 266124 100042
rect 265808 97640 265860 97646
rect 265808 97582 265860 97588
rect 265900 97096 265952 97102
rect 265900 97038 265952 97044
rect 265624 96824 265676 96830
rect 265624 96766 265676 96772
rect 264980 96756 265032 96762
rect 264980 96698 265032 96704
rect 264888 92472 264940 92478
rect 264888 92414 264940 92420
rect 264704 88120 264756 88126
rect 264704 88062 264756 88068
rect 264520 82408 264572 82414
rect 264520 82350 264572 82356
rect 265912 12170 265940 97038
rect 265992 96960 266044 96966
rect 266096 96948 266124 100014
rect 266188 97102 266216 100028
rect 266176 97096 266228 97102
rect 266176 97038 266228 97044
rect 266096 96920 266308 96948
rect 265992 96902 266044 96908
rect 266004 89622 266032 96902
rect 266176 96824 266228 96830
rect 266176 96766 266228 96772
rect 266084 96756 266136 96762
rect 266084 96698 266136 96704
rect 265992 89616 266044 89622
rect 265992 89558 266044 89564
rect 266096 12306 266124 96698
rect 266084 12300 266136 12306
rect 266084 12242 266136 12248
rect 266188 12238 266216 96766
rect 266280 92274 266308 96920
rect 266464 96830 266492 100028
rect 266648 96898 266676 100028
rect 266832 96966 266860 100028
rect 267030 100014 267136 100042
rect 267004 97028 267056 97034
rect 267004 96970 267056 96976
rect 266820 96960 266872 96966
rect 266820 96902 266872 96908
rect 266636 96892 266688 96898
rect 266636 96834 266688 96840
rect 266452 96824 266504 96830
rect 266452 96766 266504 96772
rect 267016 92342 267044 96970
rect 267108 96948 267136 100014
rect 267200 97102 267228 100028
rect 267398 100014 267504 100042
rect 267280 97776 267332 97782
rect 267280 97718 267332 97724
rect 267292 97238 267320 97718
rect 267280 97232 267332 97238
rect 267280 97174 267332 97180
rect 267188 97096 267240 97102
rect 267188 97038 267240 97044
rect 267372 96960 267424 96966
rect 267108 96920 267320 96948
rect 267188 96824 267240 96830
rect 267188 96766 267240 96772
rect 267004 92336 267056 92342
rect 267004 92278 267056 92284
rect 266268 92268 266320 92274
rect 266268 92210 266320 92216
rect 267200 88058 267228 96766
rect 267188 88052 267240 88058
rect 267188 87994 267240 88000
rect 267292 86698 267320 96920
rect 267372 96902 267424 96908
rect 267280 86692 267332 86698
rect 267280 86634 267332 86640
rect 267004 13116 267056 13122
rect 267004 13058 267056 13064
rect 266176 12232 266228 12238
rect 266176 12174 266228 12180
rect 265900 12164 265952 12170
rect 265900 12106 265952 12112
rect 265348 5228 265400 5234
rect 265348 5170 265400 5176
rect 264244 3664 264296 3670
rect 264244 3606 264296 3612
rect 265360 480 265388 5170
rect 267016 4010 267044 13058
rect 267384 12102 267412 96902
rect 267372 12096 267424 12102
rect 267372 12038 267424 12044
rect 267476 12034 267504 100014
rect 267660 98002 267688 100028
rect 267660 97974 267780 98002
rect 267648 97708 267700 97714
rect 267648 97650 267700 97656
rect 267660 97102 267688 97650
rect 267752 97510 267780 97974
rect 267740 97504 267792 97510
rect 267740 97446 267792 97452
rect 267556 97096 267608 97102
rect 267556 97038 267608 97044
rect 267648 97096 267700 97102
rect 267648 97038 267700 97044
rect 267464 12028 267516 12034
rect 267464 11970 267516 11976
rect 267568 8022 267596 97038
rect 267844 96898 267872 100028
rect 268028 96966 268056 100028
rect 268212 97782 268240 100028
rect 268200 97776 268252 97782
rect 268200 97718 268252 97724
rect 268016 96960 268068 96966
rect 268016 96902 268068 96908
rect 267648 96892 267700 96898
rect 267648 96834 267700 96840
rect 267832 96892 267884 96898
rect 267832 96834 267884 96840
rect 267660 8090 267688 96834
rect 268396 96830 268424 100028
rect 268594 100014 268792 100042
rect 268660 96960 268712 96966
rect 268660 96902 268712 96908
rect 268568 96892 268620 96898
rect 268568 96834 268620 96840
rect 268384 96824 268436 96830
rect 268384 96766 268436 96772
rect 267648 8084 267700 8090
rect 267648 8026 267700 8032
rect 267556 8016 267608 8022
rect 267556 7958 267608 7964
rect 268580 7954 268608 96834
rect 268672 11966 268700 96902
rect 268660 11960 268712 11966
rect 268660 11902 268712 11908
rect 268764 11898 268792 100014
rect 268856 97238 268884 100028
rect 268948 100014 269054 100042
rect 268844 97232 268896 97238
rect 268844 97174 268896 97180
rect 268948 96914 268976 100014
rect 269028 97232 269080 97238
rect 269028 97174 269080 97180
rect 268856 96886 268976 96914
rect 268752 11892 268804 11898
rect 268752 11834 268804 11840
rect 268568 7948 268620 7954
rect 268568 7890 268620 7896
rect 268856 7818 268884 96886
rect 268936 96824 268988 96830
rect 268936 96766 268988 96772
rect 268948 7886 268976 96766
rect 269040 90982 269068 97174
rect 269224 96762 269252 100028
rect 269408 96830 269436 100028
rect 269592 96898 269620 100028
rect 269776 96966 269804 100028
rect 270052 97238 270080 100028
rect 270144 100014 270250 100042
rect 270040 97232 270092 97238
rect 270040 97174 270092 97180
rect 269764 96960 269816 96966
rect 270144 96914 270172 100014
rect 269764 96902 269816 96908
rect 269580 96892 269632 96898
rect 269580 96834 269632 96840
rect 269960 96886 270172 96914
rect 270224 96960 270276 96966
rect 270224 96902 270276 96908
rect 269396 96824 269448 96830
rect 269396 96766 269448 96772
rect 269212 96756 269264 96762
rect 269212 96698 269264 96704
rect 269028 90976 269080 90982
rect 269028 90918 269080 90924
rect 268936 7880 268988 7886
rect 268936 7822 268988 7828
rect 268844 7812 268896 7818
rect 268844 7754 268896 7760
rect 269960 7682 269988 96886
rect 270040 96824 270092 96830
rect 270040 96766 270092 96772
rect 270052 86834 270080 96766
rect 270132 96756 270184 96762
rect 270132 96698 270184 96704
rect 270040 86828 270092 86834
rect 270040 86770 270092 86776
rect 270144 11830 270172 96698
rect 270132 11824 270184 11830
rect 270132 11766 270184 11772
rect 270236 11762 270264 96902
rect 270316 96892 270368 96898
rect 270316 96834 270368 96840
rect 270224 11756 270276 11762
rect 270224 11698 270276 11704
rect 270328 7750 270356 96834
rect 270420 93566 270448 100028
rect 270604 97714 270632 100028
rect 270788 98394 270816 100028
rect 270776 98388 270828 98394
rect 270776 98330 270828 98336
rect 270972 98326 271000 100028
rect 270960 98320 271012 98326
rect 270960 98262 271012 98268
rect 270592 97708 270644 97714
rect 270592 97650 270644 97656
rect 271052 97300 271104 97306
rect 271052 97242 271104 97248
rect 271064 93854 271092 97242
rect 271144 97232 271196 97238
rect 271144 97174 271196 97180
rect 271156 96778 271184 97174
rect 271248 96966 271276 100028
rect 271432 99210 271460 100028
rect 271630 100014 271736 100042
rect 271420 99204 271472 99210
rect 271420 99146 271472 99152
rect 271328 97436 271380 97442
rect 271328 97378 271380 97384
rect 271236 96960 271288 96966
rect 271236 96902 271288 96908
rect 271156 96750 271276 96778
rect 271064 93826 271184 93854
rect 270408 93560 270460 93566
rect 270408 93502 270460 93508
rect 270316 7744 270368 7750
rect 270316 7686 270368 7692
rect 269948 7676 270000 7682
rect 269948 7618 270000 7624
rect 268844 5024 268896 5030
rect 268844 4966 268896 4972
rect 266728 4004 266780 4010
rect 266728 3946 266780 3952
rect 267004 4004 267056 4010
rect 267004 3946 267056 3952
rect 266740 3670 266768 3946
rect 267740 3936 267792 3942
rect 267740 3878 267792 3884
rect 266728 3664 266780 3670
rect 266728 3606 266780 3612
rect 266544 3596 266596 3602
rect 266544 3538 266596 3544
rect 266556 480 266584 3538
rect 267752 480 267780 3878
rect 268856 480 268884 4966
rect 271156 3534 271184 93826
rect 271248 5030 271276 96750
rect 271340 85270 271368 97378
rect 271708 89554 271736 100014
rect 271800 97050 271828 100028
rect 271800 97022 271920 97050
rect 271788 96960 271840 96966
rect 271788 96902 271840 96908
rect 271696 89548 271748 89554
rect 271696 89490 271748 89496
rect 271328 85264 271380 85270
rect 271328 85206 271380 85212
rect 271800 82278 271828 96902
rect 271892 96762 271920 97022
rect 271984 96898 272012 100028
rect 271972 96892 272024 96898
rect 271972 96834 272024 96840
rect 272168 96830 272196 100028
rect 272444 97306 272472 100028
rect 272432 97300 272484 97306
rect 272432 97242 272484 97248
rect 272628 96966 272656 100028
rect 272708 97912 272760 97918
rect 272708 97854 272760 97860
rect 272720 97646 272748 97854
rect 272708 97640 272760 97646
rect 272708 97582 272760 97588
rect 272616 96960 272668 96966
rect 272616 96902 272668 96908
rect 272156 96824 272208 96830
rect 272156 96766 272208 96772
rect 271880 96756 271932 96762
rect 271880 96698 271932 96704
rect 272812 86630 272840 100028
rect 272996 97714 273024 100028
rect 273088 100014 273194 100042
rect 272984 97708 273036 97714
rect 272984 97650 273036 97656
rect 272892 96960 272944 96966
rect 273088 96914 273116 100014
rect 273260 97504 273312 97510
rect 273260 97446 273312 97452
rect 273272 96966 273300 97446
rect 272892 96902 272944 96908
rect 272904 92206 272932 96902
rect 272996 96886 273116 96914
rect 273260 96960 273312 96966
rect 273260 96902 273312 96908
rect 273168 96892 273220 96898
rect 272892 92200 272944 92206
rect 272892 92142 272944 92148
rect 272996 92138 273024 96886
rect 273168 96834 273220 96840
rect 273076 96824 273128 96830
rect 273076 96766 273128 96772
rect 272984 92132 273036 92138
rect 272984 92074 273036 92080
rect 273088 87990 273116 96766
rect 273180 93498 273208 96834
rect 273364 96762 273392 100028
rect 273352 96756 273404 96762
rect 273352 96698 273404 96704
rect 273640 96694 273668 100028
rect 273824 99142 273852 100028
rect 274022 100014 274128 100042
rect 273812 99136 273864 99142
rect 273812 99078 273864 99084
rect 274100 96914 274128 100014
rect 274192 97238 274220 100028
rect 274180 97232 274232 97238
rect 274180 97174 274232 97180
rect 274100 96886 274220 96914
rect 274088 96824 274140 96830
rect 274088 96766 274140 96772
rect 273628 96688 273680 96694
rect 273628 96630 273680 96636
rect 273168 93492 273220 93498
rect 273168 93434 273220 93440
rect 273076 87984 273128 87990
rect 273076 87926 273128 87932
rect 272800 86624 272852 86630
rect 272800 86566 272852 86572
rect 273904 83496 273956 83502
rect 273904 83438 273956 83444
rect 271788 82272 271840 82278
rect 271788 82214 271840 82220
rect 271236 5024 271288 5030
rect 271236 4966 271288 4972
rect 273916 4010 273944 83438
rect 274100 7614 274128 96766
rect 274192 87922 274220 96886
rect 274376 96830 274404 100028
rect 274468 100014 274574 100042
rect 274364 96824 274416 96830
rect 274364 96766 274416 96772
rect 274468 96642 274496 100014
rect 274548 97232 274600 97238
rect 274548 97174 274600 97180
rect 274284 96614 274496 96642
rect 274180 87916 274232 87922
rect 274180 87858 274232 87864
rect 274284 86562 274312 96614
rect 274364 96552 274416 96558
rect 274560 96506 274588 97174
rect 274640 96756 274692 96762
rect 274640 96698 274692 96704
rect 274364 96494 274416 96500
rect 274272 86556 274324 86562
rect 274272 86498 274324 86504
rect 274376 83774 274404 96494
rect 274468 96478 274588 96506
rect 274364 83768 274416 83774
rect 274364 83710 274416 83716
rect 274468 80782 274496 96478
rect 274652 96370 274680 96698
rect 274836 96694 274864 100028
rect 275020 99074 275048 100028
rect 275218 100014 275324 100042
rect 275008 99068 275060 99074
rect 275008 99010 275060 99016
rect 275296 96914 275324 100014
rect 275388 97782 275416 100028
rect 275376 97776 275428 97782
rect 275376 97718 275428 97724
rect 275572 97238 275600 100028
rect 275560 97232 275612 97238
rect 275560 97174 275612 97180
rect 275296 96886 275692 96914
rect 275560 96756 275612 96762
rect 275560 96698 275612 96704
rect 274824 96688 274876 96694
rect 274824 96630 274876 96636
rect 274560 96342 274680 96370
rect 274560 91050 274588 96342
rect 274548 91044 274600 91050
rect 274548 90986 274600 90992
rect 275284 82136 275336 82142
rect 275284 82078 275336 82084
rect 274456 80776 274508 80782
rect 274456 80718 274508 80724
rect 274088 7608 274140 7614
rect 274088 7550 274140 7556
rect 271236 4004 271288 4010
rect 271236 3946 271288 3952
rect 273904 4004 273956 4010
rect 273904 3946 273956 3952
rect 270040 3528 270092 3534
rect 270040 3470 270092 3476
rect 271144 3528 271196 3534
rect 271144 3470 271196 3476
rect 270052 480 270080 3470
rect 271248 480 271276 3946
rect 273628 3596 273680 3602
rect 273628 3538 273680 3544
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 272444 480 272472 3402
rect 273640 480 273668 3538
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 274836 480 274864 3470
rect 275296 2922 275324 82078
rect 275572 80850 275600 96698
rect 275664 89486 275692 96886
rect 275652 89480 275704 89486
rect 275652 89422 275704 89428
rect 275756 86494 275784 100028
rect 275848 100014 275954 100042
rect 275848 96762 275876 100014
rect 276020 97844 276072 97850
rect 276020 97786 276072 97792
rect 276032 97238 276060 97786
rect 275928 97232 275980 97238
rect 275928 97174 275980 97180
rect 276020 97232 276072 97238
rect 276020 97174 276072 97180
rect 275836 96756 275888 96762
rect 275836 96698 275888 96704
rect 275836 96552 275888 96558
rect 275836 96494 275888 96500
rect 275744 86488 275796 86494
rect 275744 86430 275796 86436
rect 275848 82346 275876 96494
rect 275940 93430 275968 97174
rect 276216 96762 276244 100028
rect 276204 96756 276256 96762
rect 276204 96698 276256 96704
rect 276400 96694 276428 100028
rect 276584 97442 276612 100028
rect 276782 100014 276888 100042
rect 276966 100014 277072 100042
rect 276572 97436 276624 97442
rect 276572 97378 276624 97384
rect 276664 97368 276716 97374
rect 276664 97310 276716 97316
rect 276756 97368 276808 97374
rect 276756 97310 276808 97316
rect 276388 96688 276440 96694
rect 276388 96630 276440 96636
rect 275928 93424 275980 93430
rect 275928 93366 275980 93372
rect 276676 83910 276704 97310
rect 276768 93854 276796 97310
rect 276860 96914 276888 100014
rect 277044 97050 277072 100014
rect 277136 97374 277164 100028
rect 277412 98938 277440 100028
rect 277400 98932 277452 98938
rect 277400 98874 277452 98880
rect 277308 97640 277360 97646
rect 277308 97582 277360 97588
rect 277124 97368 277176 97374
rect 277124 97310 277176 97316
rect 277044 97022 277164 97050
rect 276860 96886 277072 96914
rect 276768 93826 276980 93854
rect 276664 83904 276716 83910
rect 276664 83846 276716 83852
rect 275836 82340 275888 82346
rect 275836 82282 275888 82288
rect 275560 80844 275612 80850
rect 275560 80786 275612 80792
rect 276020 4956 276072 4962
rect 276020 4898 276072 4904
rect 275284 2916 275336 2922
rect 275284 2858 275336 2864
rect 276032 480 276060 4898
rect 276952 3534 276980 93826
rect 277044 92002 277072 96886
rect 277032 91996 277084 92002
rect 277032 91938 277084 91944
rect 277136 13394 277164 97022
rect 277320 96898 277348 97582
rect 277308 96892 277360 96898
rect 277308 96834 277360 96840
rect 277596 96762 277624 100028
rect 277780 97646 277808 100028
rect 277768 97640 277820 97646
rect 277768 97582 277820 97588
rect 277964 96830 277992 100028
rect 278162 100014 278268 100042
rect 278136 97844 278188 97850
rect 278136 97786 278188 97792
rect 278148 96898 278176 97786
rect 278136 96892 278188 96898
rect 278136 96834 278188 96840
rect 277952 96824 278004 96830
rect 277952 96766 278004 96772
rect 277308 96756 277360 96762
rect 277308 96698 277360 96704
rect 277584 96756 277636 96762
rect 277584 96698 277636 96704
rect 277216 96688 277268 96694
rect 277216 96630 277268 96636
rect 277228 13462 277256 96630
rect 277320 92070 277348 96698
rect 278240 93854 278268 100014
rect 278332 96898 278360 100028
rect 278424 100014 278622 100042
rect 278320 96892 278372 96898
rect 278320 96834 278372 96840
rect 278240 93826 278360 93854
rect 277308 92064 277360 92070
rect 277308 92006 277360 92012
rect 277216 13456 277268 13462
rect 277216 13398 277268 13404
rect 277124 13388 277176 13394
rect 277124 13330 277176 13336
rect 278332 13258 278360 93826
rect 278424 90846 278452 100014
rect 278504 96892 278556 96898
rect 278504 96834 278556 96840
rect 278412 90840 278464 90846
rect 278412 90782 278464 90788
rect 278516 82142 278544 96834
rect 278792 96830 278820 100028
rect 278976 97510 279004 100028
rect 279160 98870 279188 100028
rect 279148 98864 279200 98870
rect 279148 98806 279200 98812
rect 278964 97504 279016 97510
rect 278964 97446 279016 97452
rect 279344 96898 279372 100028
rect 279332 96892 279384 96898
rect 279332 96834 279384 96840
rect 278688 96824 278740 96830
rect 278688 96766 278740 96772
rect 278780 96824 278832 96830
rect 278780 96766 278832 96772
rect 278596 96756 278648 96762
rect 278596 96698 278648 96704
rect 278504 82136 278556 82142
rect 278504 82078 278556 82084
rect 278608 13326 278636 96698
rect 278700 91934 278728 96766
rect 279528 96762 279556 100028
rect 279712 100014 279818 100042
rect 279896 100014 280002 100042
rect 279516 96756 279568 96762
rect 279516 96698 279568 96704
rect 279712 95130 279740 100014
rect 279896 96914 279924 100014
rect 280172 97345 280200 100028
rect 280158 97336 280214 97345
rect 280158 97271 280214 97280
rect 279804 96886 279924 96914
rect 279976 96892 280028 96898
rect 279700 95124 279752 95130
rect 279700 95066 279752 95072
rect 278688 91928 278740 91934
rect 278688 91870 278740 91876
rect 279804 85202 279832 96886
rect 279976 96834 280028 96840
rect 279884 96824 279936 96830
rect 279884 96766 279936 96772
rect 279896 91866 279924 96766
rect 279884 91860 279936 91866
rect 279884 91802 279936 91808
rect 279988 86426 280016 96834
rect 280356 96830 280384 100028
rect 280540 96898 280568 100028
rect 280738 100014 280936 100042
rect 280528 96892 280580 96898
rect 280528 96834 280580 96840
rect 280344 96824 280396 96830
rect 280344 96766 280396 96772
rect 280908 93854 280936 100014
rect 281000 96014 281028 100028
rect 281198 100014 281304 100042
rect 281080 97300 281132 97306
rect 281080 97242 281132 97248
rect 280988 96008 281040 96014
rect 280988 95950 281040 95956
rect 280908 93826 281028 93854
rect 279976 86420 280028 86426
rect 279976 86362 280028 86368
rect 279792 85196 279844 85202
rect 279792 85138 279844 85144
rect 278596 13320 278648 13326
rect 278596 13262 278648 13268
rect 278320 13252 278372 13258
rect 278320 13194 278372 13200
rect 280712 8968 280764 8974
rect 280712 8910 280764 8916
rect 278320 4004 278372 4010
rect 278320 3946 278372 3952
rect 277124 3868 277176 3874
rect 277124 3810 277176 3816
rect 276940 3528 276992 3534
rect 276940 3470 276992 3476
rect 277136 480 277164 3810
rect 278332 480 278360 3946
rect 279516 2916 279568 2922
rect 279516 2858 279568 2864
rect 279528 480 279556 2858
rect 280724 480 280752 8910
rect 281000 3398 281028 93826
rect 281092 13122 281120 97242
rect 281276 96914 281304 100014
rect 281368 97306 281396 100028
rect 281356 97300 281408 97306
rect 281356 97242 281408 97248
rect 281172 96892 281224 96898
rect 281276 96886 281396 96914
rect 281172 96834 281224 96840
rect 281184 13190 281212 96834
rect 281264 96824 281316 96830
rect 281264 96766 281316 96772
rect 281172 13184 281224 13190
rect 281172 13126 281224 13132
rect 281080 13116 281132 13122
rect 281080 13058 281132 13064
rect 281276 9042 281304 96766
rect 281264 9036 281316 9042
rect 281264 8978 281316 8984
rect 281368 8974 281396 96886
rect 281552 96218 281580 100028
rect 281736 96898 281764 100028
rect 281724 96892 281776 96898
rect 281724 96834 281776 96840
rect 281540 96212 281592 96218
rect 281540 96154 281592 96160
rect 281920 85134 281948 100028
rect 282104 100014 282210 100042
rect 282000 97640 282052 97646
rect 281998 97608 282000 97617
rect 282052 97608 282054 97617
rect 281998 97543 282054 97552
rect 282000 97504 282052 97510
rect 282000 97446 282052 97452
rect 282012 97306 282040 97446
rect 282000 97300 282052 97306
rect 282000 97242 282052 97248
rect 282104 96286 282132 100014
rect 282184 97776 282236 97782
rect 282184 97718 282236 97724
rect 282196 97510 282224 97718
rect 282276 97708 282328 97714
rect 282276 97650 282328 97656
rect 282184 97504 282236 97510
rect 282184 97446 282236 97452
rect 282288 97374 282316 97650
rect 282276 97368 282328 97374
rect 282276 97310 282328 97316
rect 282380 96830 282408 100028
rect 282472 100014 282578 100042
rect 282762 100014 282868 100042
rect 282368 96824 282420 96830
rect 282368 96766 282420 96772
rect 282092 96280 282144 96286
rect 282092 96222 282144 96228
rect 282184 95940 282236 95946
rect 282184 95882 282236 95888
rect 281908 85128 281960 85134
rect 281908 85070 281960 85076
rect 281540 14476 281592 14482
rect 281540 14418 281592 14424
rect 281356 8968 281408 8974
rect 281356 8910 281408 8916
rect 280988 3392 281040 3398
rect 280988 3334 281040 3340
rect 281552 490 281580 14418
rect 282196 3466 282224 95882
rect 282472 19990 282500 100014
rect 282736 97776 282788 97782
rect 282736 97718 282788 97724
rect 282644 96892 282696 96898
rect 282644 96834 282696 96840
rect 282552 96824 282604 96830
rect 282552 96766 282604 96772
rect 282564 90710 282592 96766
rect 282656 90778 282684 96834
rect 282748 96694 282776 97718
rect 282736 96688 282788 96694
rect 282736 96630 282788 96636
rect 282840 96354 282868 100014
rect 282932 98802 282960 100028
rect 282920 98796 282972 98802
rect 282920 98738 282972 98744
rect 283116 96694 283144 100028
rect 283104 96688 283156 96694
rect 283104 96630 283156 96636
rect 282828 96348 282880 96354
rect 282828 96290 282880 96296
rect 283392 96150 283420 100028
rect 283576 96830 283604 100028
rect 283760 96898 283788 100028
rect 283852 100014 283958 100042
rect 284036 100014 284142 100042
rect 283748 96892 283800 96898
rect 283748 96834 283800 96840
rect 283564 96824 283616 96830
rect 283852 96778 283880 100014
rect 284036 96914 284064 100014
rect 283564 96766 283616 96772
rect 283760 96750 283880 96778
rect 283944 96886 284064 96914
rect 284312 96898 284340 100028
rect 284116 96892 284168 96898
rect 283760 96490 283788 96750
rect 283840 96688 283892 96694
rect 283840 96630 283892 96636
rect 283748 96484 283800 96490
rect 283748 96426 283800 96432
rect 283380 96144 283432 96150
rect 283380 96086 283432 96092
rect 282644 90772 282696 90778
rect 282644 90714 282696 90720
rect 282552 90704 282604 90710
rect 282552 90646 282604 90652
rect 283852 85066 283880 96630
rect 283944 90574 283972 96886
rect 284116 96834 284168 96840
rect 284300 96892 284352 96898
rect 284300 96834 284352 96840
rect 284024 96824 284076 96830
rect 284024 96766 284076 96772
rect 284036 90642 284064 96766
rect 284024 90636 284076 90642
rect 284024 90578 284076 90584
rect 283932 90568 283984 90574
rect 283932 90510 283984 90516
rect 284128 86358 284156 96834
rect 284588 96082 284616 100028
rect 284786 100014 284892 100042
rect 284970 100014 285076 100042
rect 284864 96506 284892 100014
rect 285048 96914 285076 100014
rect 285140 97306 285168 100028
rect 285128 97300 285180 97306
rect 285128 97242 285180 97248
rect 285048 96886 285260 96914
rect 284864 96478 285168 96506
rect 285036 96416 285088 96422
rect 285036 96358 285088 96364
rect 284576 96076 284628 96082
rect 284576 96018 284628 96024
rect 284116 86352 284168 86358
rect 284116 86294 284168 86300
rect 283840 85060 283892 85066
rect 283840 85002 283892 85008
rect 284300 80708 284352 80714
rect 284300 80650 284352 80656
rect 282460 19984 282512 19990
rect 282460 19926 282512 19932
rect 282184 3460 282236 3466
rect 282184 3402 282236 3408
rect 283104 3460 283156 3466
rect 283104 3402 283156 3408
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 3402
rect 284312 480 284340 80650
rect 285048 24138 285076 96358
rect 285140 90506 285168 96478
rect 285128 90500 285180 90506
rect 285128 90442 285180 90448
rect 285036 24132 285088 24138
rect 285036 24074 285088 24080
rect 285232 4962 285260 96886
rect 285324 89418 285352 100028
rect 285416 100014 285522 100042
rect 285416 96422 285444 100014
rect 285588 97300 285640 97306
rect 285588 97242 285640 97248
rect 285496 96892 285548 96898
rect 285496 96834 285548 96840
rect 285404 96416 285456 96422
rect 285404 96358 285456 96364
rect 285312 89412 285364 89418
rect 285312 89354 285364 89360
rect 285508 84998 285536 96834
rect 285600 96558 285628 97242
rect 285588 96552 285640 96558
rect 285588 96494 285640 96500
rect 285784 96014 285812 100028
rect 285862 97608 285918 97617
rect 285862 97543 285918 97552
rect 285876 97374 285904 97543
rect 285864 97368 285916 97374
rect 285864 97310 285916 97316
rect 285968 96898 285996 100028
rect 286166 100014 286272 100042
rect 285956 96892 286008 96898
rect 285956 96834 286008 96840
rect 285864 96280 285916 96286
rect 285864 96222 285916 96228
rect 285772 96008 285824 96014
rect 285772 95950 285824 95956
rect 285876 95946 285904 96222
rect 285864 95940 285916 95946
rect 285864 95882 285916 95888
rect 285680 94580 285732 94586
rect 285680 94522 285732 94528
rect 285496 84992 285548 84998
rect 285496 84934 285548 84940
rect 285220 4956 285272 4962
rect 285220 4898 285272 4904
rect 285692 3482 285720 94522
rect 286244 93854 286272 100014
rect 286336 94858 286364 100028
rect 286520 96830 286548 100028
rect 286612 100014 286718 100042
rect 286508 96824 286560 96830
rect 286508 96766 286560 96772
rect 286324 94852 286376 94858
rect 286324 94794 286376 94800
rect 286244 93826 286548 93854
rect 286520 83706 286548 93826
rect 286508 83700 286560 83706
rect 286508 83642 286560 83648
rect 286612 26926 286640 100014
rect 286692 96892 286744 96898
rect 286692 96834 286744 96840
rect 286704 90438 286732 96834
rect 286784 96824 286836 96830
rect 286784 96766 286836 96772
rect 286692 90432 286744 90438
rect 286692 90374 286744 90380
rect 286796 89350 286824 96766
rect 286980 95198 287008 100028
rect 287164 96830 287192 100028
rect 287152 96824 287204 96830
rect 287152 96766 287204 96772
rect 287348 96694 287376 100028
rect 287336 96688 287388 96694
rect 287336 96630 287388 96636
rect 287532 95470 287560 100028
rect 287716 96762 287744 100028
rect 287914 100014 288020 100042
rect 287796 96824 287848 96830
rect 287796 96766 287848 96772
rect 287704 96756 287756 96762
rect 287704 96698 287756 96704
rect 287520 95464 287572 95470
rect 287520 95406 287572 95412
rect 286968 95192 287020 95198
rect 286968 95134 287020 95140
rect 287808 91798 287836 96766
rect 287888 96688 287940 96694
rect 287888 96630 287940 96636
rect 287796 91792 287848 91798
rect 287796 91734 287848 91740
rect 286784 89344 286836 89350
rect 286784 89286 286836 89292
rect 287060 89004 287112 89010
rect 287060 88946 287112 88952
rect 286600 26920 286652 26926
rect 286600 26862 286652 26868
rect 285416 3454 285720 3482
rect 285416 480 285444 3454
rect 287072 2802 287100 88946
rect 287900 83638 287928 96630
rect 287888 83632 287940 83638
rect 287888 83574 287940 83580
rect 287992 18630 288020 100014
rect 288072 96756 288124 96762
rect 288072 96698 288124 96704
rect 288084 89282 288112 96698
rect 288176 94790 288204 100028
rect 288268 100014 288374 100042
rect 288164 94784 288216 94790
rect 288164 94726 288216 94732
rect 288072 89276 288124 89282
rect 288072 89218 288124 89224
rect 288268 89214 288296 100014
rect 288544 96762 288572 100028
rect 288532 96756 288584 96762
rect 288532 96698 288584 96704
rect 288728 94722 288756 100028
rect 288926 100014 289032 100042
rect 289110 100014 289308 100042
rect 289004 96914 289032 100014
rect 289280 97050 289308 100014
rect 289372 98258 289400 100028
rect 289464 100014 289570 100042
rect 289360 98252 289412 98258
rect 289360 98194 289412 98200
rect 289280 97022 289400 97050
rect 289004 96886 289308 96914
rect 289176 96824 289228 96830
rect 289176 96766 289228 96772
rect 288716 94716 288768 94722
rect 288716 94658 288768 94664
rect 288256 89208 288308 89214
rect 288256 89150 288308 89156
rect 289188 60042 289216 96766
rect 289280 90914 289308 96886
rect 289268 90908 289320 90914
rect 289268 90850 289320 90856
rect 289176 60036 289228 60042
rect 289176 59978 289228 59984
rect 287980 18624 288032 18630
rect 287980 18566 288032 18572
rect 287796 6724 287848 6730
rect 287796 6666 287848 6672
rect 286980 2774 287100 2802
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 2774
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 6666
rect 289372 4894 289400 97022
rect 289464 89146 289492 100014
rect 289636 98252 289688 98258
rect 289636 98194 289688 98200
rect 289544 96756 289596 96762
rect 289544 96698 289596 96704
rect 289452 89140 289504 89146
rect 289452 89082 289504 89088
rect 289556 84930 289584 96698
rect 289648 94926 289676 98194
rect 289740 96830 289768 100028
rect 289728 96824 289780 96830
rect 289728 96766 289780 96772
rect 289924 95985 289952 100028
rect 290108 99006 290136 100028
rect 290306 100014 290504 100042
rect 290096 99000 290148 99006
rect 290096 98942 290148 98948
rect 289910 95976 289966 95985
rect 289910 95911 289966 95920
rect 289636 94920 289688 94926
rect 289636 94862 289688 94868
rect 290476 86290 290504 100014
rect 290568 94654 290596 100028
rect 290752 96830 290780 100028
rect 290844 100014 290950 100042
rect 290740 96824 290792 96830
rect 290740 96766 290792 96772
rect 290556 94648 290608 94654
rect 290556 94590 290608 94596
rect 290464 86284 290516 86290
rect 290464 86226 290516 86232
rect 289544 84924 289596 84930
rect 289544 84866 289596 84872
rect 290844 83570 290872 100014
rect 290924 96824 290976 96830
rect 290924 96766 290976 96772
rect 290936 89078 290964 96766
rect 291120 94994 291148 100028
rect 291304 96830 291332 100028
rect 291292 96824 291344 96830
rect 291292 96766 291344 96772
rect 291488 96762 291516 100028
rect 291476 96756 291528 96762
rect 291476 96698 291528 96704
rect 291108 94988 291160 94994
rect 291108 94930 291160 94936
rect 291764 94586 291792 100028
rect 291856 100014 291962 100042
rect 292040 100014 292146 100042
rect 291856 96694 291884 100014
rect 291936 96824 291988 96830
rect 291936 96766 291988 96772
rect 291844 96688 291896 96694
rect 291844 96630 291896 96636
rect 291752 94580 291804 94586
rect 291752 94522 291804 94528
rect 291948 90370 291976 96766
rect 291936 90364 291988 90370
rect 291936 90306 291988 90312
rect 290924 89072 290976 89078
rect 290924 89014 290976 89020
rect 290832 83564 290884 83570
rect 290832 83506 290884 83512
rect 292040 21418 292068 100014
rect 292212 96824 292264 96830
rect 292212 96766 292264 96772
rect 292316 96778 292344 100028
rect 292500 96830 292528 100028
rect 292488 96824 292540 96830
rect 292120 96756 292172 96762
rect 292120 96698 292172 96704
rect 292028 21412 292080 21418
rect 292028 21354 292080 21360
rect 292132 6186 292160 96698
rect 292224 87718 292252 96766
rect 292316 96750 292436 96778
rect 292488 96766 292540 96772
rect 292304 96688 292356 96694
rect 292304 96630 292356 96636
rect 292316 87786 292344 96630
rect 292408 95062 292436 96750
rect 292396 95056 292448 95062
rect 292396 94998 292448 95004
rect 292684 94110 292712 100028
rect 292960 98734 292988 100028
rect 292948 98728 293000 98734
rect 292948 98670 293000 98676
rect 293144 95849 293172 100028
rect 293342 100014 293448 100042
rect 293130 95840 293186 95849
rect 293130 95775 293186 95784
rect 293420 94518 293448 100014
rect 293512 98666 293540 100028
rect 293710 100014 293816 100042
rect 293500 98660 293552 98666
rect 293500 98602 293552 98608
rect 293788 96778 293816 100014
rect 293512 96750 293816 96778
rect 293224 94512 293276 94518
rect 293224 94454 293276 94460
rect 293408 94512 293460 94518
rect 293408 94454 293460 94460
rect 292672 94104 292724 94110
rect 292672 94046 292724 94052
rect 292304 87780 292356 87786
rect 292304 87722 292356 87728
rect 292212 87712 292264 87718
rect 292212 87654 292264 87660
rect 291384 6180 291436 6186
rect 291384 6122 291436 6128
rect 292120 6180 292172 6186
rect 292120 6122 292172 6128
rect 290188 5160 290240 5166
rect 290188 5102 290240 5108
rect 288992 4888 289044 4894
rect 288992 4830 289044 4836
rect 289360 4888 289412 4894
rect 289360 4830 289412 4836
rect 289004 480 289032 4830
rect 290200 480 290228 5102
rect 291396 480 291424 6122
rect 292580 4820 292632 4826
rect 292580 4762 292632 4768
rect 292592 480 292620 4762
rect 293236 3602 293264 94454
rect 293512 93362 293540 96750
rect 293880 94602 293908 100028
rect 294156 96694 294184 100028
rect 294354 100014 294460 100042
rect 294432 96830 294460 100014
rect 294420 96824 294472 96830
rect 294420 96766 294472 96772
rect 294524 96762 294552 100028
rect 294512 96756 294564 96762
rect 294512 96698 294564 96704
rect 294144 96688 294196 96694
rect 294144 96630 294196 96636
rect 293604 94574 293908 94602
rect 293500 93356 293552 93362
rect 293500 93298 293552 93304
rect 293604 83502 293632 94574
rect 293776 94512 293828 94518
rect 293776 94454 293828 94460
rect 293684 94104 293736 94110
rect 293684 94046 293736 94052
rect 293696 87854 293724 94046
rect 293684 87848 293736 87854
rect 293684 87790 293736 87796
rect 293788 84862 293816 94454
rect 294708 93294 294736 100028
rect 294906 100014 295012 100042
rect 295090 100014 295196 100042
rect 294984 99374 295012 100014
rect 294984 99346 295104 99374
rect 294972 96756 295024 96762
rect 294972 96698 295024 96704
rect 294788 96688 294840 96694
rect 294788 96630 294840 96636
rect 294880 96688 294932 96694
rect 294880 96630 294932 96636
rect 294696 93288 294748 93294
rect 294696 93230 294748 93236
rect 293776 84856 293828 84862
rect 293776 84798 293828 84804
rect 293592 83496 293644 83502
rect 293592 83438 293644 83444
rect 293684 5092 293736 5098
rect 293684 5034 293736 5040
rect 293224 3596 293276 3602
rect 293224 3538 293276 3544
rect 293696 480 293724 5034
rect 294800 4826 294828 96630
rect 294892 14618 294920 96630
rect 294984 14686 295012 96698
rect 294972 14680 295024 14686
rect 294972 14622 295024 14628
rect 294880 14612 294932 14618
rect 294880 14554 294932 14560
rect 295076 10470 295104 99346
rect 295168 96694 295196 100014
rect 295248 96824 295300 96830
rect 295248 96766 295300 96772
rect 295156 96688 295208 96694
rect 295156 96630 295208 96636
rect 295260 89714 295288 96766
rect 295352 94518 295380 100028
rect 295536 96830 295564 100028
rect 295524 96824 295576 96830
rect 295524 96766 295576 96772
rect 295720 96694 295748 100028
rect 295918 100014 296024 100042
rect 295708 96688 295760 96694
rect 295708 96630 295760 96636
rect 295340 94512 295392 94518
rect 295340 94454 295392 94460
rect 295996 93226 296024 100014
rect 296088 96762 296116 100028
rect 296076 96756 296128 96762
rect 296076 96698 296128 96704
rect 296168 96688 296220 96694
rect 296168 96630 296220 96636
rect 295984 93220 296036 93226
rect 295984 93162 296036 93168
rect 295168 89686 295288 89714
rect 295168 10538 295196 89686
rect 296180 82210 296208 96630
rect 296168 82204 296220 82210
rect 296168 82146 296220 82152
rect 295984 82136 296036 82142
rect 295984 82078 296036 82084
rect 295156 10532 295208 10538
rect 295156 10474 295208 10480
rect 295064 10464 295116 10470
rect 295064 10406 295116 10412
rect 294788 4820 294840 4826
rect 294788 4762 294840 4768
rect 295996 3602 296024 82078
rect 296272 22778 296300 100028
rect 296444 96824 296496 96830
rect 296444 96766 296496 96772
rect 296352 96756 296404 96762
rect 296352 96698 296404 96704
rect 296364 89010 296392 96698
rect 296352 89004 296404 89010
rect 296352 88946 296404 88952
rect 296456 87650 296484 96766
rect 296548 93158 296576 100028
rect 296732 96830 296760 100028
rect 296930 100014 297036 100042
rect 296720 96824 296772 96830
rect 296720 96766 296772 96772
rect 297008 96762 297036 100014
rect 296996 96756 297048 96762
rect 296996 96698 297048 96704
rect 297100 96665 297128 100028
rect 297284 96694 297312 100028
rect 297482 100014 297680 100042
rect 297272 96688 297324 96694
rect 297086 96656 297142 96665
rect 297272 96630 297324 96636
rect 297086 96591 297142 96600
rect 297364 95940 297416 95946
rect 297364 95882 297416 95888
rect 297376 95470 297404 95882
rect 297364 95464 297416 95470
rect 297364 95406 297416 95412
rect 296536 93152 296588 93158
rect 296536 93094 296588 93100
rect 297652 89714 297680 100014
rect 297744 97209 297772 100028
rect 297928 97481 297956 100028
rect 298112 99374 298140 100028
rect 298296 99414 298324 100028
rect 298284 99408 298336 99414
rect 298112 99346 298232 99374
rect 298284 99350 298336 99356
rect 298480 99346 298508 100028
rect 298664 99618 298692 100028
rect 298940 99754 298968 100028
rect 298928 99748 298980 99754
rect 298928 99690 298980 99696
rect 299124 99686 299152 100028
rect 299112 99680 299164 99686
rect 299112 99622 299164 99628
rect 298652 99612 298704 99618
rect 298652 99554 298704 99560
rect 297914 97472 297970 97481
rect 297914 97407 297970 97416
rect 297730 97200 297786 97209
rect 297730 97135 297786 97144
rect 298008 97164 298060 97170
rect 298008 97106 298060 97112
rect 298020 96762 298048 97106
rect 298204 96830 298232 99346
rect 298468 99340 298520 99346
rect 298468 99282 298520 99288
rect 299308 99278 299336 100028
rect 299492 99550 299520 100028
rect 299480 99544 299532 99550
rect 299480 99486 299532 99492
rect 299676 99414 299704 100028
rect 299860 99482 299888 100028
rect 299848 99476 299900 99482
rect 299848 99418 299900 99424
rect 299664 99408 299716 99414
rect 299664 99350 299716 99356
rect 301516 99346 301544 122062
rect 302516 120080 302568 120086
rect 302516 120022 302568 120028
rect 302528 119921 302556 120022
rect 302514 119912 302570 119921
rect 302514 119847 302570 119856
rect 302608 117292 302660 117298
rect 302608 117234 302660 117240
rect 302620 116929 302648 117234
rect 302606 116920 302662 116929
rect 302606 116855 302662 116864
rect 302516 111784 302568 111790
rect 302516 111726 302568 111732
rect 302528 110673 302556 111726
rect 302514 110664 302570 110673
rect 302514 110599 302570 110608
rect 302792 108996 302844 109002
rect 302792 108938 302844 108944
rect 302804 107681 302832 108938
rect 302790 107672 302846 107681
rect 302790 107607 302846 107616
rect 302896 104553 302924 123422
rect 302988 113801 303016 123490
rect 302974 113792 303030 113801
rect 302974 113727 303030 113736
rect 302882 104544 302938 104553
rect 302882 104479 302938 104488
rect 302792 102128 302844 102134
rect 302792 102070 302844 102076
rect 302804 101561 302832 102070
rect 302790 101552 302846 101561
rect 302790 101487 302846 101496
rect 305748 99346 305776 193802
rect 307680 152930 307708 251194
rect 307668 152924 307720 152930
rect 307668 152866 307720 152872
rect 309796 122602 309824 302194
rect 312544 301504 312596 301510
rect 312544 301446 312596 301452
rect 311164 300212 311216 300218
rect 311164 300154 311216 300160
rect 309784 122596 309836 122602
rect 309784 122538 309836 122544
rect 301504 99340 301556 99346
rect 301504 99282 301556 99288
rect 305736 99340 305788 99346
rect 305736 99282 305788 99288
rect 299296 99272 299348 99278
rect 299296 99214 299348 99220
rect 302884 97164 302936 97170
rect 302884 97106 302936 97112
rect 300124 97028 300176 97034
rect 300124 96970 300176 96976
rect 298836 96960 298888 96966
rect 298836 96902 298888 96908
rect 298100 96824 298152 96830
rect 298100 96766 298152 96772
rect 298192 96824 298244 96830
rect 298192 96766 298244 96772
rect 297824 96756 297876 96762
rect 297824 96698 297876 96704
rect 298008 96756 298060 96762
rect 298008 96698 298060 96704
rect 297652 89686 297772 89714
rect 296444 87644 296496 87650
rect 296444 87586 296496 87592
rect 296260 22772 296312 22778
rect 296260 22714 296312 22720
rect 297744 14482 297772 89686
rect 297836 14550 297864 96698
rect 297916 96688 297968 96694
rect 298112 96642 298140 96766
rect 297916 96630 297968 96636
rect 297824 14544 297876 14550
rect 297824 14486 297876 14492
rect 297732 14476 297784 14482
rect 297732 14418 297784 14424
rect 297928 10334 297956 96630
rect 298020 96614 298140 96642
rect 298742 96656 298798 96665
rect 298020 10402 298048 96614
rect 298742 96591 298798 96600
rect 298192 95600 298244 95606
rect 298192 95542 298244 95548
rect 298100 16108 298152 16114
rect 298100 16050 298152 16056
rect 298008 10396 298060 10402
rect 298008 10338 298060 10344
rect 297916 10328 297968 10334
rect 297916 10270 297968 10276
rect 297272 6248 297324 6254
rect 297272 6190 297324 6196
rect 296076 4004 296128 4010
rect 296076 3946 296128 3952
rect 294880 3596 294932 3602
rect 294880 3538 294932 3544
rect 295984 3596 296036 3602
rect 295984 3538 296036 3544
rect 294892 480 294920 3538
rect 296088 480 296116 3946
rect 297284 480 297312 6190
rect 298112 490 298140 16050
rect 298204 4010 298232 95542
rect 298756 80714 298784 96591
rect 298848 82482 298876 96902
rect 299480 95532 299532 95538
rect 299480 95474 299532 95480
rect 298836 82476 298888 82482
rect 298836 82418 298888 82424
rect 298744 80708 298796 80714
rect 298744 80650 298796 80656
rect 298192 4004 298244 4010
rect 298192 3946 298244 3952
rect 299492 3482 299520 95474
rect 299572 10940 299624 10946
rect 299572 10882 299624 10888
rect 299584 3874 299612 10882
rect 300136 9110 300164 96970
rect 302240 95736 302292 95742
rect 302240 95678 302292 95684
rect 302252 16574 302280 95678
rect 302252 16546 302832 16574
rect 301504 16040 301556 16046
rect 301504 15982 301556 15988
rect 300124 9104 300176 9110
rect 300124 9046 300176 9052
rect 299572 3868 299624 3874
rect 299572 3810 299624 3816
rect 300768 3868 300820 3874
rect 300768 3810 300820 3816
rect 299492 3454 299704 3482
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3454
rect 300780 480 300808 3810
rect 301516 490 301544 15982
rect 302804 3482 302832 16546
rect 302896 5098 302924 97106
rect 307024 96892 307076 96898
rect 307024 96834 307076 96840
rect 304356 96824 304408 96830
rect 304356 96766 304408 96772
rect 304264 96756 304316 96762
rect 304264 96698 304316 96704
rect 303896 10872 303948 10878
rect 303896 10814 303948 10820
rect 302884 5092 302936 5098
rect 302884 5034 302936 5040
rect 302804 3454 303200 3482
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 3454
rect 303908 490 303936 10814
rect 304276 3942 304304 96698
rect 304368 82142 304396 96766
rect 306380 95668 306432 95674
rect 306380 95610 306432 95616
rect 304356 82136 304408 82142
rect 304356 82078 304408 82084
rect 304264 3936 304316 3942
rect 304264 3878 304316 3884
rect 305552 3732 305604 3738
rect 305552 3674 305604 3680
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3674
rect 306392 490 306420 95610
rect 307036 6254 307064 96834
rect 309140 95804 309192 95810
rect 309140 95746 309192 95752
rect 309152 16574 309180 95746
rect 311176 86970 311204 300154
rect 312556 245614 312584 301446
rect 318064 301436 318116 301442
rect 318064 301378 318116 301384
rect 313924 301368 313976 301374
rect 313924 301310 313976 301316
rect 313188 258732 313240 258738
rect 313188 258674 313240 258680
rect 313200 258126 313228 258674
rect 313188 258120 313240 258126
rect 313188 258062 313240 258068
rect 312544 245608 312596 245614
rect 312544 245550 312596 245556
rect 313200 152862 313228 258062
rect 313188 152856 313240 152862
rect 313188 152798 313240 152804
rect 312544 95872 312596 95878
rect 312544 95814 312596 95820
rect 311256 88800 311308 88806
rect 311256 88742 311308 88748
rect 311164 86964 311216 86970
rect 311164 86906 311216 86912
rect 309152 16546 309824 16574
rect 307760 15972 307812 15978
rect 307760 15914 307812 15920
rect 307024 6248 307076 6254
rect 307024 6190 307076 6196
rect 307772 3398 307800 15914
rect 307944 10804 307996 10810
rect 307944 10746 307996 10752
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 10746
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 309796 490 309824 16546
rect 311164 10736 311216 10742
rect 311164 10678 311216 10684
rect 311176 3210 311204 10678
rect 311268 3398 311296 88742
rect 311256 3392 311308 3398
rect 311256 3334 311308 3340
rect 311176 3182 311480 3210
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 3182
rect 312556 2990 312584 95814
rect 313280 94240 313332 94246
rect 313280 94182 313332 94188
rect 313292 16574 313320 94182
rect 313936 33114 313964 301310
rect 316684 300144 316736 300150
rect 316684 300086 316736 300092
rect 316040 94308 316092 94314
rect 316040 94250 316092 94256
rect 313924 33108 313976 33114
rect 313924 33050 313976 33056
rect 313292 16546 313872 16574
rect 312636 3392 312688 3398
rect 312636 3334 312688 3340
rect 312544 2984 312596 2990
rect 312544 2926 312596 2932
rect 312648 480 312676 3334
rect 313844 480 313872 16546
rect 316052 3398 316080 94250
rect 316696 73166 316724 300086
rect 318076 113150 318104 301378
rect 320824 295384 320876 295390
rect 320824 295326 320876 295332
rect 320836 122874 320864 295326
rect 320824 122868 320876 122874
rect 320824 122810 320876 122816
rect 318064 113144 318116 113150
rect 318064 113086 318116 113092
rect 322216 99754 322244 337418
rect 322204 99748 322256 99754
rect 322204 99690 322256 99696
rect 323596 99686 323624 482394
rect 331232 330546 331260 702986
rect 348804 700942 348832 703520
rect 348792 700936 348844 700942
rect 348792 700878 348844 700884
rect 364996 699718 365024 703520
rect 397472 699718 397500 703520
rect 413664 700738 413692 703520
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 359464 699712 359516 699718
rect 359464 699654 359516 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 331220 330540 331272 330546
rect 331220 330482 331272 330488
rect 359476 305930 359504 699654
rect 371238 585712 371294 585721
rect 371238 585647 371294 585656
rect 371252 578218 371280 585647
rect 371700 585404 371752 585410
rect 371700 585346 371752 585352
rect 371712 585177 371740 585346
rect 371698 585168 371754 585177
rect 371698 585103 371754 585112
rect 371422 584624 371478 584633
rect 371422 584559 371478 584568
rect 371330 581904 371386 581913
rect 371330 581839 371386 581848
rect 371344 581058 371372 581839
rect 371332 581052 371384 581058
rect 371332 580994 371384 581000
rect 371436 579714 371464 584559
rect 371712 582298 371740 585103
rect 371792 584384 371844 584390
rect 371792 584326 371844 584332
rect 371804 582457 371832 584326
rect 371790 582448 371846 582457
rect 371790 582383 371846 582392
rect 372158 582448 372214 582457
rect 372158 582383 372214 582392
rect 371712 582270 371832 582298
rect 371606 581360 371662 581369
rect 371606 581295 371662 581304
rect 371620 581126 371648 581295
rect 371608 581120 371660 581126
rect 371608 581062 371660 581068
rect 371698 580816 371754 580825
rect 371698 580751 371754 580760
rect 371514 580272 371570 580281
rect 371514 580207 371570 580216
rect 371528 579834 371556 580207
rect 371516 579828 371568 579834
rect 371516 579770 371568 579776
rect 371608 579760 371660 579766
rect 371606 579728 371608 579737
rect 371660 579728 371662 579737
rect 371436 579686 371556 579714
rect 371330 578640 371386 578649
rect 371330 578575 371386 578584
rect 371344 578338 371372 578575
rect 371332 578332 371384 578338
rect 371332 578274 371384 578280
rect 371252 578190 371372 578218
rect 371240 578128 371292 578134
rect 371240 578070 371292 578076
rect 369858 569256 369914 569265
rect 369858 569191 369914 569200
rect 369306 568712 369362 568721
rect 369306 568647 369362 568656
rect 369320 567194 369348 568647
rect 369044 567166 369348 567194
rect 360212 556022 360962 556050
rect 360212 514754 360240 556022
rect 362880 553489 362908 556036
rect 364904 553489 364932 556036
rect 366928 554198 366956 556036
rect 366916 554192 366968 554198
rect 366916 554134 366968 554140
rect 362866 553480 362922 553489
rect 362866 553415 362922 553424
rect 364890 553480 364946 553489
rect 364890 553415 364946 553424
rect 368952 551954 368980 556036
rect 368940 551948 368992 551954
rect 368940 551890 368992 551896
rect 369044 514754 369072 567166
rect 369306 566536 369362 566545
rect 369306 566471 369362 566480
rect 369320 557534 369348 566471
rect 369136 557506 369348 557534
rect 369136 517002 369164 557506
rect 369308 551948 369360 551954
rect 369308 551890 369360 551896
rect 369124 516996 369176 517002
rect 369124 516938 369176 516944
rect 360212 514726 360608 514754
rect 369044 514726 369164 514754
rect 360580 484106 360608 514726
rect 369136 511834 369164 514726
rect 369124 511828 369176 511834
rect 369124 511770 369176 511776
rect 369136 507854 369164 511770
rect 369044 507826 369164 507854
rect 369044 487154 369072 507826
rect 369124 505572 369176 505578
rect 369124 505514 369176 505520
rect 369136 491366 369164 505514
rect 369320 494054 369348 551890
rect 369492 516996 369544 517002
rect 369492 516938 369544 516944
rect 369398 511864 369454 511873
rect 369398 511799 369400 511808
rect 369452 511799 369454 511808
rect 369400 511770 369452 511776
rect 369504 507521 369532 516938
rect 369872 512961 369900 569191
rect 369950 567216 370006 567225
rect 369950 567151 370006 567160
rect 369858 512952 369914 512961
rect 369858 512887 369914 512896
rect 369490 507512 369546 507521
rect 369490 507447 369546 507456
rect 369504 505578 369532 507447
rect 369492 505572 369544 505578
rect 369492 505514 369544 505520
rect 369228 494026 369348 494054
rect 369124 491360 369176 491366
rect 369124 491302 369176 491308
rect 369044 487126 369164 487154
rect 369136 484906 369164 487126
rect 369124 484900 369176 484906
rect 369124 484842 369176 484848
rect 369228 484786 369256 494026
rect 369308 491360 369360 491366
rect 369308 491302 369360 491308
rect 368966 484758 369256 484786
rect 369124 484696 369176 484702
rect 369124 484638 369176 484644
rect 365166 484120 365222 484129
rect 360580 484078 360962 484106
rect 360856 482798 360884 484078
rect 362880 483002 362908 484092
rect 364918 484078 365166 484106
rect 365166 484055 365222 484064
rect 362868 482996 362920 483002
rect 362868 482938 362920 482944
rect 360844 482792 360896 482798
rect 360844 482734 360896 482740
rect 360856 412026 360884 482734
rect 362880 482225 362908 482938
rect 366928 482458 366956 484092
rect 366916 482452 366968 482458
rect 366916 482394 366968 482400
rect 362866 482216 362922 482225
rect 362866 482151 362922 482160
rect 369136 476114 369164 484638
rect 369228 482866 369256 484758
rect 369216 482860 369268 482866
rect 369216 482802 369268 482808
rect 369044 476086 369164 476114
rect 369044 426442 369072 476086
rect 369320 470594 369348 491302
rect 369766 488200 369822 488209
rect 369766 488135 369822 488144
rect 369780 488102 369808 488135
rect 369400 488096 369452 488102
rect 369400 488038 369452 488044
rect 369768 488096 369820 488102
rect 369768 488038 369820 488044
rect 369136 470566 369348 470594
rect 369136 441614 369164 470566
rect 369136 441586 369348 441614
rect 369044 426426 369164 426442
rect 369044 426420 369176 426426
rect 369044 426414 369124 426420
rect 369124 426362 369176 426368
rect 369320 423201 369348 441586
rect 369306 423192 369362 423201
rect 369306 423127 369362 423136
rect 369306 421016 369362 421025
rect 369306 420951 369362 420960
rect 369320 412634 369348 420951
rect 369412 413953 369440 488038
rect 369768 482860 369820 482866
rect 369768 482802 369820 482808
rect 369492 426420 369544 426426
rect 369492 426362 369544 426368
rect 369504 425241 369532 426362
rect 369490 425232 369546 425241
rect 369490 425167 369546 425176
rect 369398 413944 369454 413953
rect 369398 413879 369454 413888
rect 369228 412606 369348 412634
rect 369124 412072 369176 412078
rect 362774 412040 362830 412049
rect 360580 411998 360962 412026
rect 360580 393314 360608 411998
rect 365166 412040 365222 412049
rect 362830 411998 362894 412026
rect 364918 411998 365166 412026
rect 362774 411975 362830 411984
rect 368966 412020 369124 412026
rect 368966 412014 369176 412020
rect 365166 411975 365222 411984
rect 366928 409222 366956 412012
rect 368966 411998 369164 412014
rect 366916 409216 366968 409222
rect 366916 409158 366968 409164
rect 360212 393286 360608 393314
rect 360212 369854 360240 393286
rect 360212 369826 360608 369854
rect 360580 340082 360608 369826
rect 362498 340504 362554 340513
rect 365166 340504 365222 340513
rect 362554 340462 362894 340490
rect 364918 340462 365166 340490
rect 362498 340439 362554 340448
rect 365166 340439 365222 340448
rect 369044 340082 369072 411998
rect 369228 383654 369256 412606
rect 369780 412078 369808 482802
rect 369872 425921 369900 512887
rect 369964 509425 369992 567151
rect 370134 564224 370190 564233
rect 370134 564159 370190 564168
rect 369950 509416 370006 509425
rect 369950 509351 370006 509360
rect 369858 425912 369914 425921
rect 369858 425847 369914 425856
rect 369964 423609 369992 509351
rect 370044 505504 370096 505510
rect 370044 505446 370096 505452
rect 370056 504937 370084 505446
rect 370042 504928 370098 504937
rect 370042 504863 370098 504872
rect 369950 423600 370006 423609
rect 369950 423535 370006 423544
rect 370056 421705 370084 504863
rect 370148 501945 370176 564159
rect 370226 562048 370282 562057
rect 370226 561983 370282 561992
rect 370134 501936 370190 501945
rect 370134 501871 370190 501880
rect 370042 421696 370098 421705
rect 370042 421631 370098 421640
rect 369950 417752 370006 417761
rect 369950 417687 370006 417696
rect 369768 412072 369820 412078
rect 369768 412014 369820 412020
rect 369858 411632 369914 411641
rect 369858 411567 369914 411576
rect 369228 383626 369348 383654
rect 369124 363588 369176 363594
rect 369124 363530 369176 363536
rect 360580 340054 360962 340082
rect 368966 340068 369072 340082
rect 360580 335354 360608 340054
rect 366928 337482 366956 340068
rect 368952 340054 369072 340068
rect 368952 339250 368980 340054
rect 368940 339244 368992 339250
rect 368940 339186 368992 339192
rect 366916 337476 366968 337482
rect 366916 337418 366968 337424
rect 360212 335326 360608 335354
rect 359464 305924 359516 305930
rect 359464 305866 359516 305872
rect 347688 296200 347740 296206
rect 347688 296142 347740 296148
rect 347700 258738 347728 296142
rect 358084 296064 358136 296070
rect 358084 296006 358136 296012
rect 353944 282940 353996 282946
rect 353944 282882 353996 282888
rect 353956 266218 353984 282882
rect 356704 278792 356756 278798
rect 356704 278734 356756 278740
rect 353944 266212 353996 266218
rect 353944 266154 353996 266160
rect 356716 266121 356744 278734
rect 356702 266112 356758 266121
rect 356702 266047 356758 266056
rect 358096 264926 358124 296006
rect 359464 295860 359516 295866
rect 359464 295802 359516 295808
rect 358176 276072 358228 276078
rect 358176 276014 358228 276020
rect 358188 266257 358216 276014
rect 358174 266248 358230 266257
rect 358174 266183 358230 266192
rect 358084 264920 358136 264926
rect 358084 264862 358136 264868
rect 359476 262206 359504 295802
rect 360212 287054 360240 335326
rect 360212 287026 360608 287054
rect 360580 273290 360608 287026
rect 369136 283506 369164 363530
rect 369320 359825 369348 383626
rect 369306 359816 369362 359825
rect 369306 359751 369362 359760
rect 369320 342254 369348 359751
rect 369768 359168 369820 359174
rect 369768 359110 369820 359116
rect 369780 358873 369808 359110
rect 369766 358864 369822 358873
rect 369766 358799 369822 358808
rect 369780 357814 369808 358799
rect 369768 357808 369820 357814
rect 369768 357750 369820 357756
rect 369228 342226 369348 342254
rect 369228 283626 369256 342226
rect 369872 340921 369900 411567
rect 369964 353569 369992 417687
rect 370056 360913 370084 421631
rect 370148 420209 370176 501871
rect 370240 497321 370268 561983
rect 370318 561504 370374 561513
rect 370318 561439 370374 561448
rect 370226 497312 370282 497321
rect 370226 497247 370282 497256
rect 370134 420200 370190 420209
rect 370134 420135 370190 420144
rect 370042 360904 370098 360913
rect 370042 360839 370098 360848
rect 369950 353560 370006 353569
rect 369950 353495 370006 353504
rect 369858 340912 369914 340921
rect 369858 340847 369914 340856
rect 369308 339244 369360 339250
rect 369308 339186 369360 339192
rect 369216 283620 369268 283626
rect 369216 283562 369268 283568
rect 369136 283478 369256 283506
rect 369124 283348 369176 283354
rect 369124 283290 369176 283296
rect 360568 273284 360620 273290
rect 369136 273254 369164 283290
rect 369228 280906 369256 283478
rect 369216 280900 369268 280906
rect 369216 280842 369268 280848
rect 369320 277394 369348 339186
rect 369398 297528 369454 297537
rect 369398 297463 369400 297472
rect 369452 297463 369454 297472
rect 369400 297434 369452 297440
rect 369860 297424 369912 297430
rect 369858 297392 369860 297401
rect 369912 297392 369914 297401
rect 369858 297327 369914 297336
rect 369400 296200 369452 296206
rect 369400 296142 369452 296148
rect 369412 295905 369440 296142
rect 369398 295896 369454 295905
rect 369398 295831 369454 295840
rect 369858 295896 369914 295905
rect 369858 295831 369860 295840
rect 369912 295831 369914 295840
rect 369860 295802 369912 295808
rect 369490 291952 369546 291961
rect 369490 291887 369546 291896
rect 369398 283384 369454 283393
rect 369398 283319 369400 283328
rect 369452 283319 369454 283328
rect 369400 283290 369452 283296
rect 369400 280900 369452 280906
rect 369400 280842 369452 280848
rect 369412 280809 369440 280842
rect 369398 280800 369454 280809
rect 369398 280735 369454 280744
rect 360568 273226 360620 273232
rect 369044 273226 369164 273254
rect 369228 277366 369348 277394
rect 360580 268138 360608 273226
rect 369044 270494 369072 273226
rect 369044 270466 369164 270494
rect 369136 268258 369164 270466
rect 369124 268252 369176 268258
rect 369124 268194 369176 268200
rect 369228 268138 369256 277366
rect 360580 268124 360962 268138
rect 368966 268124 369256 268138
rect 360580 268110 360976 268124
rect 360948 265742 360976 268110
rect 362880 266354 362908 268124
rect 362868 266348 362920 266354
rect 362868 266290 362920 266296
rect 362880 266257 362908 266290
rect 364904 266286 364932 268124
rect 364892 266280 364944 266286
rect 362866 266248 362922 266257
rect 364892 266222 364944 266228
rect 362866 266183 362922 266192
rect 364904 265849 364932 266222
rect 366928 266150 366956 268124
rect 368952 268110 369256 268124
rect 368952 266218 368980 268110
rect 369032 268048 369084 268054
rect 369032 267990 369084 267996
rect 368940 266212 368992 266218
rect 368940 266154 368992 266160
rect 366916 266144 366968 266150
rect 366916 266086 366968 266092
rect 364890 265840 364946 265849
rect 364890 265775 364946 265784
rect 360200 265736 360252 265742
rect 360200 265678 360252 265684
rect 360936 265736 360988 265742
rect 360936 265678 360988 265684
rect 359464 262200 359516 262206
rect 359464 262142 359516 262148
rect 357348 260160 357400 260166
rect 357348 260102 357400 260108
rect 347688 258732 347740 258738
rect 347688 258674 347740 258680
rect 357360 256018 357388 260102
rect 357348 256012 357400 256018
rect 357348 255954 357400 255960
rect 357360 255338 357388 255954
rect 357348 255332 357400 255338
rect 357348 255274 357400 255280
rect 340328 246356 340380 246362
rect 340328 246298 340380 246304
rect 340340 245682 340368 246298
rect 340328 245676 340380 245682
rect 340328 245618 340380 245624
rect 340788 245676 340840 245682
rect 340788 245618 340840 245624
rect 340800 152726 340828 245618
rect 342904 242208 342956 242214
rect 342904 242150 342956 242156
rect 340880 224392 340932 224398
rect 340880 224334 340932 224340
rect 340892 223922 340920 224334
rect 340880 223916 340932 223922
rect 340880 223858 340932 223864
rect 342168 223916 342220 223922
rect 342168 223858 342220 223864
rect 342180 153066 342208 223858
rect 342916 209098 342944 242150
rect 351920 225072 351972 225078
rect 351920 225014 351972 225020
rect 345664 225004 345716 225010
rect 345664 224946 345716 224952
rect 345676 219434 345704 224946
rect 351932 222154 351960 225014
rect 351920 222148 351972 222154
rect 351920 222090 351972 222096
rect 345664 219428 345716 219434
rect 345664 219370 345716 219376
rect 352564 215960 352616 215966
rect 352564 215902 352616 215908
rect 342904 209092 342956 209098
rect 342904 209034 342956 209040
rect 346308 199436 346360 199442
rect 346308 199378 346360 199384
rect 346320 195362 346348 199378
rect 346308 195356 346360 195362
rect 346308 195298 346360 195304
rect 352576 189786 352604 215902
rect 352564 189780 352616 189786
rect 352564 189722 352616 189728
rect 357256 175296 357308 175302
rect 357256 175238 357308 175244
rect 342168 153060 342220 153066
rect 342168 153002 342220 153008
rect 357268 152794 357296 175238
rect 357360 152998 357388 255274
rect 360212 224954 360240 265678
rect 367834 225720 367890 225729
rect 367834 225655 367836 225664
rect 367888 225655 367890 225664
rect 367836 225626 367888 225632
rect 360212 224926 360608 224954
rect 358084 224324 358136 224330
rect 358084 224266 358136 224272
rect 358096 175302 358124 224266
rect 360580 196738 360608 224926
rect 369044 204254 369072 267990
rect 369124 266212 369176 266218
rect 369124 266154 369176 266160
rect 369136 218054 369164 266154
rect 369412 224954 369440 280735
rect 369504 264246 369532 291887
rect 369950 287872 370006 287881
rect 369950 287807 370006 287816
rect 369858 284472 369914 284481
rect 369858 284407 369914 284416
rect 369676 283620 369728 283626
rect 369676 283562 369728 283568
rect 369688 277545 369716 283562
rect 369674 277536 369730 277545
rect 369674 277471 369730 277480
rect 369492 264240 369544 264246
rect 369492 264182 369544 264188
rect 369412 224926 369532 224954
rect 369400 224324 369452 224330
rect 369400 224266 369452 224272
rect 369412 224233 369440 224266
rect 369398 224224 369454 224233
rect 369398 224159 369454 224168
rect 369504 223689 369532 224926
rect 369490 223680 369546 223689
rect 369490 223615 369546 223624
rect 369136 218026 369348 218054
rect 369044 204226 369256 204254
rect 369124 197396 369176 197402
rect 369124 197338 369176 197344
rect 360580 196710 360962 196738
rect 359464 194472 359516 194478
rect 359464 194414 359516 194420
rect 358084 175296 358136 175302
rect 358084 175238 358136 175244
rect 359004 153332 359056 153338
rect 359004 153274 359056 153280
rect 357348 152992 357400 152998
rect 357348 152934 357400 152940
rect 357256 152788 357308 152794
rect 357256 152730 357308 152736
rect 340788 152720 340840 152726
rect 340788 152662 340840 152668
rect 359016 151774 359044 153274
rect 359004 151768 359056 151774
rect 359004 151710 359056 151716
rect 323584 99680 323636 99686
rect 323584 99622 323636 99628
rect 359476 99618 359504 194414
rect 360580 180794 360608 196710
rect 365166 196480 365222 196489
rect 364918 196438 365166 196466
rect 365166 196415 365222 196424
rect 369136 196058 369164 197338
rect 362880 194585 362908 196044
rect 362866 194576 362922 194585
rect 362866 194511 362922 194520
rect 366928 194478 366956 196044
rect 368966 196030 369164 196058
rect 366916 194472 366968 194478
rect 366916 194414 366968 194420
rect 360212 180766 360608 180794
rect 359648 154012 359700 154018
rect 359648 153954 359700 153960
rect 359556 151904 359608 151910
rect 359556 151846 359608 151852
rect 359568 142118 359596 151846
rect 359660 144906 359688 153954
rect 359648 144900 359700 144906
rect 359648 144842 359700 144848
rect 359556 142112 359608 142118
rect 359556 142054 359608 142060
rect 360212 132494 360240 180766
rect 368388 176656 368440 176662
rect 368388 176598 368440 176604
rect 368400 154562 368428 176598
rect 369032 164212 369084 164218
rect 369032 164154 369084 164160
rect 369044 162926 369072 164154
rect 369032 162920 369084 162926
rect 369032 162862 369084 162868
rect 368388 154556 368440 154562
rect 368388 154498 368440 154504
rect 368400 154018 368428 154498
rect 368388 154012 368440 154018
rect 368388 153954 368440 153960
rect 369044 134994 369072 162862
rect 369136 135250 369164 196030
rect 369228 191826 369256 204226
rect 369320 197402 369348 218026
rect 369308 197396 369360 197402
rect 369308 197338 369360 197344
rect 369872 197266 369900 284407
rect 369964 268462 369992 287807
rect 370056 278089 370084 360839
rect 370148 357921 370176 420135
rect 370240 418033 370268 497247
rect 370332 496233 370360 561439
rect 370410 558240 370466 558249
rect 370410 558175 370466 558184
rect 370318 496224 370374 496233
rect 370318 496159 370374 496168
rect 370424 489394 370452 558175
rect 370504 556844 370556 556850
rect 370504 556786 370556 556792
rect 370516 556209 370544 556786
rect 370502 556200 370558 556209
rect 370502 556135 370558 556144
rect 370412 489388 370464 489394
rect 370412 489330 370464 489336
rect 370424 489297 370452 489330
rect 370410 489288 370466 489297
rect 370410 489223 370466 489232
rect 370516 484673 370544 556135
rect 370964 511216 371016 511222
rect 370962 511184 370964 511193
rect 371016 511184 371018 511193
rect 370962 511119 371018 511128
rect 370962 510096 371018 510105
rect 370962 510031 370964 510040
rect 371016 510031 371018 510040
rect 370964 510002 371016 510008
rect 370962 506560 371018 506569
rect 370962 506495 370964 506504
rect 371016 506495 371018 506504
rect 370964 506466 371016 506472
rect 370962 504248 371018 504257
rect 370962 504183 370964 504192
rect 371016 504183 371018 504192
rect 370964 504154 371016 504160
rect 370964 503192 371016 503198
rect 370962 503160 370964 503169
rect 371016 503160 371018 503169
rect 370962 503095 371018 503104
rect 370964 499656 371016 499662
rect 370962 499624 370964 499633
rect 371016 499624 371018 499633
rect 370962 499559 371018 499568
rect 370962 498536 371018 498545
rect 370962 498471 370964 498480
rect 371016 498471 371018 498480
rect 370964 498442 371016 498448
rect 370686 496224 370742 496233
rect 370686 496159 370742 496168
rect 370700 492538 370728 496159
rect 370962 495000 371018 495009
rect 370962 494935 371018 494944
rect 370976 494834 371004 494935
rect 370964 494828 371016 494834
rect 370964 494770 371016 494776
rect 370964 494012 371016 494018
rect 370964 493954 371016 493960
rect 370976 493921 371004 493954
rect 370962 493912 371018 493921
rect 370962 493847 371018 493856
rect 370780 493332 370832 493338
rect 370780 493274 370832 493280
rect 370792 492697 370820 493274
rect 370778 492688 370834 492697
rect 370778 492623 370834 492632
rect 370700 492510 370820 492538
rect 370688 489388 370740 489394
rect 370688 489330 370740 489336
rect 370502 484664 370558 484673
rect 370502 484599 370558 484608
rect 370410 422512 370466 422521
rect 370410 422447 370466 422456
rect 370226 418024 370282 418033
rect 370226 417959 370282 417968
rect 370226 414216 370282 414225
rect 370226 414151 370282 414160
rect 370134 357912 370190 357921
rect 370134 357847 370190 357856
rect 370136 357808 370188 357814
rect 370136 357750 370188 357756
rect 370042 278080 370098 278089
rect 370042 278015 370098 278024
rect 370148 277394 370176 357750
rect 370240 345273 370268 414151
rect 370320 367532 370372 367538
rect 370320 367474 370372 367480
rect 370332 367169 370360 367474
rect 370318 367160 370374 367169
rect 370318 367095 370374 367104
rect 370332 363594 370360 367095
rect 370424 363769 370452 422447
rect 370516 412185 370544 484599
rect 370700 414225 370728 489330
rect 370792 422294 370820 492510
rect 370872 492380 370924 492386
rect 370872 492322 370924 492328
rect 370884 491609 370912 492322
rect 370870 491600 370926 491609
rect 370870 491535 370926 491544
rect 370962 490376 371018 490385
rect 370962 490311 370964 490320
rect 371016 490311 371018 490320
rect 370964 490282 371016 490288
rect 370962 485752 371018 485761
rect 370962 485687 371018 485696
rect 370976 485314 371004 485687
rect 370964 485308 371016 485314
rect 370964 485250 371016 485256
rect 371148 482928 371200 482934
rect 371146 482896 371148 482905
rect 371200 482896 371202 482905
rect 371146 482831 371202 482840
rect 371252 441674 371280 578070
rect 371344 441833 371372 578190
rect 371422 577552 371478 577561
rect 371422 577487 371478 577496
rect 371436 577046 371464 577487
rect 371424 577040 371476 577046
rect 371424 576982 371476 576988
rect 371528 576854 371556 579686
rect 371712 579698 371740 580751
rect 371606 579663 371662 579672
rect 371700 579692 371752 579698
rect 371700 579634 371752 579640
rect 371698 579184 371754 579193
rect 371698 579119 371754 579128
rect 371712 578270 371740 579119
rect 371700 578264 371752 578270
rect 371700 578206 371752 578212
rect 371804 578134 371832 582270
rect 371792 578128 371844 578134
rect 371698 578096 371754 578105
rect 371792 578070 371844 578076
rect 371698 578031 371754 578040
rect 371606 577008 371662 577017
rect 371606 576943 371608 576952
rect 371660 576943 371662 576952
rect 371608 576914 371660 576920
rect 371712 576910 371740 578031
rect 371436 576826 371556 576854
rect 371700 576904 371752 576910
rect 371700 576846 371752 576852
rect 371330 441824 371386 441833
rect 371330 441759 371386 441768
rect 371160 441646 371280 441674
rect 371160 441614 371188 441646
rect 371160 441586 371280 441614
rect 371252 441153 371280 441586
rect 371238 441144 371294 441153
rect 371238 441079 371294 441088
rect 371252 440473 371280 441079
rect 371238 440464 371294 440473
rect 371238 440399 371294 440408
rect 371240 440292 371292 440298
rect 371240 440234 371292 440240
rect 371252 432290 371280 440234
rect 371344 432410 371372 441759
rect 371436 440609 371464 576826
rect 371698 576464 371754 576473
rect 371698 576399 371754 576408
rect 371608 576156 371660 576162
rect 371608 576098 371660 576104
rect 371620 575521 371648 576098
rect 371712 575550 371740 576399
rect 371882 576056 371938 576065
rect 371882 575991 371938 576000
rect 371700 575544 371752 575550
rect 371606 575512 371662 575521
rect 371528 575470 371606 575498
rect 371528 570738 371556 575470
rect 371700 575486 371752 575492
rect 371606 575447 371662 575456
rect 371790 574968 371846 574977
rect 371790 574903 371846 574912
rect 371606 571704 371662 571713
rect 371606 571639 371662 571648
rect 371620 571538 371648 571639
rect 371608 571532 371660 571538
rect 371608 571474 371660 571480
rect 371698 571160 371754 571169
rect 371698 571095 371754 571104
rect 371528 570710 371648 570738
rect 371514 570616 371570 570625
rect 371514 570551 371570 570560
rect 371528 570314 371556 570551
rect 371516 570308 371568 570314
rect 371516 570250 371568 570256
rect 371620 570194 371648 570710
rect 371528 570166 371648 570194
rect 371528 568562 371556 570166
rect 371606 570072 371662 570081
rect 371606 570007 371608 570016
rect 371660 570007 371662 570016
rect 371608 569978 371660 569984
rect 371712 569974 371740 571095
rect 371700 569968 371752 569974
rect 371700 569910 371752 569916
rect 371528 568534 371740 568562
rect 371514 568440 371570 568449
rect 371514 568375 371570 568384
rect 371528 567934 371556 568375
rect 371516 567928 371568 567934
rect 371516 567870 371568 567876
rect 371606 567896 371662 567905
rect 371606 567831 371662 567840
rect 371516 567792 371568 567798
rect 371516 567734 371568 567740
rect 371422 440600 371478 440609
rect 371422 440535 371478 440544
rect 371436 440298 371464 440535
rect 371424 440292 371476 440298
rect 371424 440234 371476 440240
rect 371528 438410 371556 567734
rect 371620 567730 371648 567831
rect 371712 567798 371740 568534
rect 371700 567792 371752 567798
rect 371700 567734 371752 567740
rect 371608 567724 371660 567730
rect 371608 567666 371660 567672
rect 371804 567610 371832 574903
rect 371436 438382 371556 438410
rect 371620 567582 371832 567610
rect 371436 432478 371464 438382
rect 371620 438274 371648 567582
rect 371896 567194 371924 575991
rect 371974 573880 372030 573889
rect 371974 573815 372030 573824
rect 371528 438246 371648 438274
rect 371712 567166 371924 567194
rect 371424 432472 371476 432478
rect 371424 432414 371476 432420
rect 371332 432404 371384 432410
rect 371332 432346 371384 432352
rect 371252 432262 371464 432290
rect 371332 432200 371384 432206
rect 371332 432142 371384 432148
rect 371238 427408 371294 427417
rect 371238 427343 371294 427352
rect 371252 426426 371280 427343
rect 371240 426420 371292 426426
rect 371240 426362 371292 426368
rect 371054 425504 371110 425513
rect 371054 425439 371110 425448
rect 371068 424726 371096 425439
rect 371238 424960 371294 424969
rect 371238 424895 371294 424904
rect 371056 424720 371108 424726
rect 371056 424662 371108 424668
rect 371146 423328 371202 423337
rect 371146 423263 371202 423272
rect 370792 422266 370912 422294
rect 370884 417489 370912 422266
rect 371160 421666 371188 423263
rect 371252 422618 371280 424895
rect 371240 422612 371292 422618
rect 371240 422554 371292 422560
rect 371148 421660 371200 421666
rect 371148 421602 371200 421608
rect 370870 417480 370926 417489
rect 370870 417415 370926 417424
rect 370686 414216 370742 414225
rect 370686 414151 370742 414160
rect 370502 412176 370558 412185
rect 370502 412111 370558 412120
rect 370594 368384 370650 368393
rect 370594 368319 370650 368328
rect 370608 367810 370636 368319
rect 370596 367804 370648 367810
rect 370596 367746 370648 367752
rect 370410 363760 370466 363769
rect 370410 363695 370466 363704
rect 370778 363760 370834 363769
rect 370778 363695 370834 363704
rect 370320 363588 370372 363594
rect 370320 363530 370372 363536
rect 370686 357912 370742 357921
rect 370686 357847 370688 357856
rect 370740 357847 370742 357856
rect 370688 357818 370740 357824
rect 370594 353288 370650 353297
rect 370594 353223 370650 353232
rect 370608 350946 370636 353223
rect 370688 351212 370740 351218
rect 370688 351154 370740 351160
rect 370700 350985 370728 351154
rect 370686 350976 370742 350985
rect 370596 350940 370648 350946
rect 370686 350911 370742 350920
rect 370596 350882 370648 350888
rect 370502 347576 370558 347585
rect 370502 347511 370558 347520
rect 370516 347206 370544 347511
rect 370504 347200 370556 347206
rect 370504 347142 370556 347148
rect 370226 345264 370282 345273
rect 370226 345199 370228 345208
rect 370280 345199 370282 345208
rect 370228 345170 370280 345176
rect 370240 345139 370268 345170
rect 370226 340640 370282 340649
rect 370226 340575 370282 340584
rect 370056 277366 370176 277394
rect 370056 277001 370084 277366
rect 370042 276992 370098 277001
rect 370042 276927 370098 276936
rect 369952 268456 370004 268462
rect 369952 268398 370004 268404
rect 369952 268320 370004 268326
rect 369952 268262 370004 268268
rect 369964 268025 369992 268262
rect 369950 268016 370006 268025
rect 369950 267951 370006 267960
rect 369860 197260 369912 197266
rect 369860 197202 369912 197208
rect 369872 196654 369900 197202
rect 369964 196897 369992 267951
rect 370056 229094 370084 276927
rect 370240 268326 370268 340575
rect 370502 295080 370558 295089
rect 370502 295015 370558 295024
rect 370410 285424 370466 285433
rect 370410 285359 370466 285368
rect 370318 278896 370374 278905
rect 370318 278831 370374 278840
rect 370228 268320 370280 268326
rect 370228 268262 370280 268268
rect 370228 266212 370280 266218
rect 370228 266154 370280 266160
rect 370240 265674 370268 266154
rect 370228 265668 370280 265674
rect 370228 265610 370280 265616
rect 370056 229066 370176 229094
rect 370148 215121 370176 229066
rect 370332 220930 370360 278831
rect 370424 250510 370452 285359
rect 370516 260166 370544 295015
rect 370594 294536 370650 294545
rect 370594 294471 370650 294480
rect 370608 267034 370636 294471
rect 370686 292904 370742 292913
rect 370686 292839 370742 292848
rect 370700 268394 370728 292839
rect 370792 278905 370820 363695
rect 370884 352209 370912 417415
rect 371238 415304 371294 415313
rect 371238 415239 371294 415248
rect 371252 414050 371280 415239
rect 371240 414044 371292 414050
rect 371240 413986 371292 413992
rect 371238 413672 371294 413681
rect 371238 413607 371294 413616
rect 371252 412146 371280 413607
rect 371240 412140 371292 412146
rect 371240 412082 371292 412088
rect 370962 369472 371018 369481
rect 370962 369407 371018 369416
rect 370976 369374 371004 369407
rect 370964 369368 371016 369374
rect 370964 369310 371016 369316
rect 371344 367198 371372 432142
rect 371436 368558 371464 432262
rect 371528 430953 371556 438246
rect 371608 438184 371660 438190
rect 371608 438126 371660 438132
rect 371620 437889 371648 438126
rect 371606 437880 371662 437889
rect 371606 437815 371662 437824
rect 371712 437442 371740 567166
rect 371790 566264 371846 566273
rect 371790 566199 371792 566208
rect 371844 566199 371846 566208
rect 371792 566170 371844 566176
rect 371792 565888 371844 565894
rect 371790 565856 371792 565865
rect 371844 565856 371846 565865
rect 371790 565791 371846 565800
rect 371790 564768 371846 564777
rect 371790 564703 371792 564712
rect 371844 564703 371846 564712
rect 371792 564674 371844 564680
rect 371790 563136 371846 563145
rect 371790 563071 371792 563080
rect 371844 563071 371846 563080
rect 371792 563042 371844 563048
rect 371790 562592 371846 562601
rect 371790 562527 371792 562536
rect 371844 562527 371846 562536
rect 371792 562498 371844 562504
rect 371790 560960 371846 560969
rect 371790 560895 371792 560904
rect 371844 560895 371846 560904
rect 371792 560866 371844 560872
rect 371790 560416 371846 560425
rect 371790 560351 371792 560360
rect 371844 560351 371846 560360
rect 371792 560322 371844 560328
rect 371882 559872 371938 559881
rect 371882 559807 371938 559816
rect 371790 559328 371846 559337
rect 371790 559263 371846 559272
rect 371804 559162 371832 559263
rect 371792 559156 371844 559162
rect 371792 559098 371844 559104
rect 371896 558958 371924 559807
rect 371884 558952 371936 558958
rect 371884 558894 371936 558900
rect 371790 558784 371846 558793
rect 371790 558719 371846 558728
rect 371804 558210 371832 558719
rect 371792 558204 371844 558210
rect 371792 558146 371844 558152
rect 371792 558068 371844 558074
rect 371792 558010 371844 558016
rect 371804 557705 371832 558010
rect 371790 557696 371846 557705
rect 371790 557631 371846 557640
rect 371790 556608 371846 556617
rect 371790 556543 371846 556552
rect 371804 556306 371832 556543
rect 371792 556300 371844 556306
rect 371792 556242 371844 556248
rect 371882 440464 371938 440473
rect 371882 440399 371938 440408
rect 371792 438932 371844 438938
rect 371792 438874 371844 438880
rect 371804 438433 371832 438874
rect 371790 438424 371846 438433
rect 371790 438359 371846 438368
rect 371700 437436 371752 437442
rect 371700 437378 371752 437384
rect 371792 437368 371844 437374
rect 371698 437336 371754 437345
rect 371608 437300 371660 437306
rect 371792 437310 371844 437316
rect 371698 437271 371754 437280
rect 371608 437242 371660 437248
rect 371620 436801 371648 437242
rect 371712 436830 371740 437271
rect 371700 436824 371752 436830
rect 371606 436792 371662 436801
rect 371700 436766 371752 436772
rect 371606 436727 371662 436736
rect 371804 436257 371832 437310
rect 371790 436248 371846 436257
rect 371790 436183 371846 436192
rect 371700 436076 371752 436082
rect 371700 436018 371752 436024
rect 371608 436008 371660 436014
rect 371608 435950 371660 435956
rect 371620 435713 371648 435950
rect 371606 435704 371662 435713
rect 371606 435639 371662 435648
rect 371712 435169 371740 436018
rect 371698 435160 371754 435169
rect 371698 435095 371754 435104
rect 371700 434716 371752 434722
rect 371700 434658 371752 434664
rect 371606 434616 371662 434625
rect 371606 434551 371608 434560
rect 371660 434551 371662 434560
rect 371608 434522 371660 434528
rect 371712 434081 371740 434658
rect 371792 434648 371844 434654
rect 371792 434590 371844 434596
rect 371698 434072 371754 434081
rect 371698 434007 371754 434016
rect 371804 433537 371832 434590
rect 371790 433528 371846 433537
rect 371790 433463 371846 433472
rect 371698 432984 371754 432993
rect 371698 432919 371754 432928
rect 371608 432676 371660 432682
rect 371608 432618 371660 432624
rect 371620 432449 371648 432618
rect 371712 432614 371740 432919
rect 371700 432608 371752 432614
rect 371700 432550 371752 432556
rect 371700 432472 371752 432478
rect 371606 432440 371662 432449
rect 371700 432414 371752 432420
rect 371606 432375 371662 432384
rect 371608 432200 371660 432206
rect 371608 432142 371660 432148
rect 371620 432041 371648 432142
rect 371606 432032 371662 432041
rect 371606 431967 371662 431976
rect 371514 430944 371570 430953
rect 371514 430879 371570 430888
rect 371424 368552 371476 368558
rect 371424 368494 371476 368500
rect 371332 367192 371384 367198
rect 371332 367134 371384 367140
rect 370964 366512 371016 366518
rect 370964 366454 371016 366460
rect 370976 366081 371004 366454
rect 370962 366072 371018 366081
rect 370962 366007 371018 366016
rect 370962 364848 371018 364857
rect 370962 364783 370964 364792
rect 371016 364783 371018 364792
rect 370964 364754 371016 364760
rect 370962 362536 371018 362545
rect 370962 362471 370964 362480
rect 371016 362471 371018 362480
rect 370964 362442 371016 362448
rect 370962 356824 371018 356833
rect 370962 356759 370964 356768
rect 371016 356759 371018 356768
rect 370964 356730 371016 356736
rect 370962 355600 371018 355609
rect 370962 355535 370964 355544
rect 371016 355535 371018 355544
rect 370964 355506 371016 355512
rect 370962 354512 371018 354521
rect 370962 354447 370964 354456
rect 371016 354447 371018 354456
rect 370964 354418 371016 354424
rect 370870 352200 370926 352209
rect 370870 352135 370872 352144
rect 370924 352135 370926 352144
rect 370872 352106 370924 352112
rect 370884 352075 370912 352106
rect 370962 349888 371018 349897
rect 370962 349823 370964 349832
rect 371016 349823 371018 349832
rect 370964 349794 371016 349800
rect 370964 348696 371016 348702
rect 370962 348664 370964 348673
rect 371016 348664 371018 348673
rect 370962 348599 371018 348608
rect 370962 346352 371018 346361
rect 370962 346287 370964 346296
rect 371016 346287 371018 346296
rect 370964 346258 371016 346264
rect 370962 344040 371018 344049
rect 370962 343975 370964 343984
rect 371016 343975 371018 343984
rect 370964 343946 371016 343952
rect 370962 342952 371018 342961
rect 370962 342887 370964 342896
rect 371016 342887 371018 342896
rect 370964 342858 371016 342864
rect 371238 298072 371294 298081
rect 371344 298042 371372 367134
rect 371436 299878 371464 368494
rect 371424 299872 371476 299878
rect 371424 299814 371476 299820
rect 371238 298007 371294 298016
rect 371332 298036 371384 298042
rect 371252 296682 371280 298007
rect 371332 297978 371384 297984
rect 371344 297809 371372 297978
rect 371330 297800 371386 297809
rect 371330 297735 371386 297744
rect 371436 296721 371464 299814
rect 371422 296712 371478 296721
rect 371240 296676 371292 296682
rect 371422 296647 371478 296656
rect 371240 296618 371292 296624
rect 371252 296206 371280 296618
rect 371240 296200 371292 296206
rect 371240 296142 371292 296148
rect 371436 296070 371464 296647
rect 371424 296064 371476 296070
rect 371424 296006 371476 296012
rect 371436 295361 371464 296006
rect 371422 295352 371478 295361
rect 371332 295316 371384 295322
rect 371422 295287 371478 295296
rect 371332 295258 371384 295264
rect 371344 294545 371372 295258
rect 371330 294536 371386 294545
rect 371330 294471 371386 294480
rect 371240 293956 371292 293962
rect 371240 293898 371292 293904
rect 371252 292913 371280 293898
rect 371332 293888 371384 293894
rect 371332 293830 371384 293836
rect 371344 293457 371372 293830
rect 371330 293448 371386 293457
rect 371330 293383 371386 293392
rect 371238 292904 371294 292913
rect 371238 292839 371294 292848
rect 371240 292528 371292 292534
rect 371240 292470 371292 292476
rect 371252 292369 371280 292470
rect 371238 292360 371294 292369
rect 371238 292295 371294 292304
rect 371332 290692 371384 290698
rect 371332 290634 371384 290640
rect 371238 289640 371294 289649
rect 371238 289575 371294 289584
rect 371252 289134 371280 289575
rect 371240 289128 371292 289134
rect 371240 289070 371292 289076
rect 371344 287609 371372 290634
rect 371330 287600 371386 287609
rect 371330 287535 371386 287544
rect 371344 287054 371372 287535
rect 371528 287065 371556 430879
rect 371620 429570 371648 431967
rect 371712 431497 371740 432414
rect 371896 431954 371924 440399
rect 371804 431926 371924 431954
rect 371698 431488 371754 431497
rect 371698 431423 371754 431432
rect 371712 430681 371740 431423
rect 371698 430672 371754 430681
rect 371698 430607 371754 430616
rect 371620 429542 371740 429570
rect 371606 427136 371662 427145
rect 371606 427071 371608 427080
rect 371660 427071 371662 427080
rect 371608 427042 371660 427048
rect 371608 426624 371660 426630
rect 371606 426592 371608 426601
rect 371660 426592 371662 426601
rect 371606 426527 371662 426536
rect 371608 426080 371660 426086
rect 371606 426048 371608 426057
rect 371660 426048 371662 426057
rect 371606 425983 371662 425992
rect 371606 423872 371662 423881
rect 371606 423807 371608 423816
rect 371660 423807 371662 423816
rect 371608 423778 371660 423784
rect 371608 423700 371660 423706
rect 371608 423642 371660 423648
rect 371068 287026 371372 287054
rect 371514 287056 371570 287065
rect 370778 278896 370834 278905
rect 370778 278831 370834 278840
rect 370688 268388 370740 268394
rect 370688 268330 370740 268336
rect 370596 267028 370648 267034
rect 370596 266970 370648 266976
rect 370504 260160 370556 260166
rect 370504 260102 370556 260108
rect 370412 250504 370464 250510
rect 370412 250446 370464 250452
rect 370412 249076 370464 249082
rect 370412 249018 370464 249024
rect 370424 248470 370452 249018
rect 370412 248464 370464 248470
rect 370412 248406 370464 248412
rect 370320 220924 370372 220930
rect 370320 220866 370372 220872
rect 370332 219745 370360 220866
rect 370318 219736 370374 219745
rect 370318 219671 370374 219680
rect 370318 218512 370374 218521
rect 370318 218447 370320 218456
rect 370372 218447 370374 218456
rect 370320 218418 370372 218424
rect 370134 215112 370190 215121
rect 370134 215047 370190 215056
rect 369950 196888 370006 196897
rect 369950 196823 370006 196832
rect 369860 196648 369912 196654
rect 369860 196590 369912 196596
rect 370320 195288 370372 195294
rect 370320 195230 370372 195236
rect 369216 191820 369268 191826
rect 369216 191762 369268 191768
rect 369400 158024 369452 158030
rect 369400 157966 369452 157972
rect 369412 155990 369440 157966
rect 369860 156664 369912 156670
rect 369860 156606 369912 156612
rect 369400 155984 369452 155990
rect 369400 155926 369452 155932
rect 369216 153196 369268 153202
rect 369216 153138 369268 153144
rect 369228 152658 369256 153138
rect 369308 152856 369360 152862
rect 369308 152798 369360 152804
rect 369216 152652 369268 152658
rect 369216 152594 369268 152600
rect 369228 146962 369256 152594
rect 369320 151745 369348 152798
rect 369306 151736 369362 151745
rect 369306 151671 369362 151680
rect 369228 146934 369348 146962
rect 369216 146872 369268 146878
rect 369216 146814 369268 146820
rect 369228 135266 369256 146814
rect 369320 136649 369348 146934
rect 369412 143857 369440 155926
rect 369676 154556 369728 154562
rect 369676 154498 369728 154504
rect 369492 152992 369544 152998
rect 369492 152934 369544 152940
rect 369504 151337 369532 152934
rect 369584 152924 369636 152930
rect 369584 152866 369636 152872
rect 369490 151328 369546 151337
rect 369490 151263 369546 151272
rect 369596 150793 369624 152866
rect 369582 150784 369638 150793
rect 369582 150719 369638 150728
rect 369398 143848 369454 143857
rect 369398 143783 369454 143792
rect 369688 142154 369716 154498
rect 369872 153270 369900 156606
rect 370136 156052 370188 156058
rect 370136 155994 370188 156000
rect 370044 153944 370096 153950
rect 370044 153886 370096 153892
rect 369860 153264 369912 153270
rect 369860 153206 369912 153212
rect 369768 151768 369820 151774
rect 369768 151710 369820 151716
rect 369780 146878 369808 151710
rect 369768 146872 369820 146878
rect 369768 146814 369820 146820
rect 369504 142126 369716 142154
rect 369306 136640 369362 136649
rect 369306 136575 369362 136584
rect 369124 135244 369176 135250
rect 369228 135238 369440 135266
rect 369124 135186 369176 135192
rect 369306 135008 369362 135017
rect 369044 134966 369306 134994
rect 369306 134943 369362 134952
rect 369124 134904 369176 134910
rect 369124 134846 369176 134852
rect 360212 132466 360608 132494
rect 360580 124794 360608 132466
rect 369136 124794 369164 134846
rect 369412 131481 369440 135238
rect 369504 132025 369532 142126
rect 369872 132433 369900 153206
rect 370056 153134 370084 153886
rect 370044 153128 370096 153134
rect 370044 153070 370096 153076
rect 370044 152584 370096 152590
rect 370044 152526 370096 152532
rect 370056 133657 370084 152526
rect 370148 139777 370176 155994
rect 370228 155236 370280 155242
rect 370228 155178 370280 155184
rect 370240 154698 370268 155178
rect 370228 154692 370280 154698
rect 370228 154634 370280 154640
rect 370240 141953 370268 154634
rect 370332 148889 370360 195230
rect 370424 149977 370452 248406
rect 371068 247722 371096 287026
rect 371514 286991 371570 287000
rect 371148 286408 371200 286414
rect 371148 286350 371200 286356
rect 371160 285977 371188 286350
rect 371528 286346 371556 286991
rect 371620 286414 371648 423642
rect 371712 296714 371740 429542
rect 371804 369578 371832 431926
rect 371882 430672 371938 430681
rect 371882 430607 371938 430616
rect 371792 369572 371844 369578
rect 371792 369514 371844 369520
rect 371804 297265 371832 369514
rect 371790 297256 371846 297265
rect 371790 297191 371846 297200
rect 371804 296818 371832 297191
rect 371792 296812 371844 296818
rect 371792 296754 371844 296760
rect 371712 296686 371832 296714
rect 371700 295248 371752 295254
rect 371700 295190 371752 295196
rect 371712 294001 371740 295190
rect 371698 293992 371754 294001
rect 371698 293927 371754 293936
rect 371700 291848 371752 291854
rect 371698 291816 371700 291825
rect 371752 291816 371754 291825
rect 371698 291751 371754 291760
rect 371698 291272 371754 291281
rect 371698 291207 371700 291216
rect 371752 291207 371754 291216
rect 371700 291178 371752 291184
rect 371698 290728 371754 290737
rect 371698 290663 371754 290672
rect 371712 290562 371740 290663
rect 371804 290578 371832 296686
rect 371896 290698 371924 430607
rect 371988 429865 372016 573815
rect 372066 573336 372122 573345
rect 372066 573271 372122 573280
rect 372080 442270 372108 573271
rect 372068 442264 372120 442270
rect 372068 442206 372120 442212
rect 371974 429856 372030 429865
rect 371974 429791 372030 429800
rect 371988 423706 372016 429791
rect 372080 429321 372108 442206
rect 372172 438938 372200 582383
rect 374000 581120 374052 581126
rect 374000 581062 374052 581068
rect 372434 574424 372490 574433
rect 372434 574359 372490 574368
rect 372250 572792 372306 572801
rect 372250 572727 372306 572736
rect 372264 556073 372292 572727
rect 372250 556064 372306 556073
rect 372250 555999 372306 556008
rect 372160 438932 372212 438938
rect 372160 438874 372212 438880
rect 372160 437436 372212 437442
rect 372160 437378 372212 437384
rect 372172 433294 372200 437378
rect 372160 433288 372212 433294
rect 372160 433230 372212 433236
rect 372172 432206 372200 433230
rect 372160 432200 372212 432206
rect 372160 432142 372212 432148
rect 372160 432064 372212 432070
rect 372160 432006 372212 432012
rect 372172 430409 372200 432006
rect 372158 430400 372214 430409
rect 372158 430335 372214 430344
rect 372066 429312 372122 429321
rect 372066 429247 372122 429256
rect 372080 429214 372108 429247
rect 372068 429208 372120 429214
rect 372068 429150 372120 429156
rect 371976 423700 372028 423706
rect 371976 423642 372028 423648
rect 372172 422294 372200 430335
rect 372264 428777 372292 555999
rect 372448 432070 372476 574359
rect 372988 567928 373040 567934
rect 372988 567870 373040 567876
rect 372526 565312 372582 565321
rect 372582 565270 372660 565298
rect 372526 565247 372582 565256
rect 372632 504218 372660 565270
rect 372710 563680 372766 563689
rect 372710 563615 372766 563624
rect 372620 504212 372672 504218
rect 372620 504154 372672 504160
rect 372526 500848 372582 500857
rect 372724 500834 372752 563615
rect 372802 557152 372858 557161
rect 372802 557087 372858 557096
rect 372582 500806 372752 500834
rect 372526 500783 372582 500792
rect 372724 500342 372752 500806
rect 372712 500336 372764 500342
rect 372712 500278 372764 500284
rect 372526 486976 372582 486985
rect 372816 486962 372844 557087
rect 372896 556300 372948 556306
rect 372896 556242 372948 556248
rect 372582 486934 372844 486962
rect 372526 486911 372582 486920
rect 372436 432064 372488 432070
rect 372436 432006 372488 432012
rect 372528 429208 372580 429214
rect 372528 429150 372580 429156
rect 372250 428768 372306 428777
rect 372250 428703 372306 428712
rect 372080 422266 372200 422294
rect 371974 422240 372030 422249
rect 371974 422175 372030 422184
rect 371988 421598 372016 422175
rect 371976 421592 372028 421598
rect 371976 421534 372028 421540
rect 371976 420776 372028 420782
rect 371974 420744 371976 420753
rect 372028 420744 372030 420753
rect 371974 420679 372030 420688
rect 371976 419144 372028 419150
rect 371974 419112 371976 419121
rect 372028 419112 372030 419121
rect 371974 419047 372030 419056
rect 371976 417444 372028 417450
rect 371976 417386 372028 417392
rect 371988 416945 372016 417386
rect 371974 416936 372030 416945
rect 371974 416871 372030 416880
rect 371976 416424 372028 416430
rect 371974 416392 371976 416401
rect 372028 416392 372030 416401
rect 371974 416327 372030 416336
rect 371974 415848 372030 415857
rect 371974 415783 372030 415792
rect 371988 415682 372016 415783
rect 371976 415676 372028 415682
rect 371976 415618 372028 415624
rect 371976 414792 372028 414798
rect 371974 414760 371976 414769
rect 372028 414760 372030 414769
rect 371974 414695 372030 414704
rect 372080 414610 372108 422266
rect 372436 419824 372488 419830
rect 372436 419766 372488 419772
rect 372448 419665 372476 419766
rect 372434 419656 372490 419665
rect 372434 419591 372490 419600
rect 372158 418568 372214 418577
rect 372158 418503 372214 418512
rect 372172 418198 372200 418503
rect 372160 418192 372212 418198
rect 372160 418134 372212 418140
rect 371988 414582 372108 414610
rect 371884 290692 371936 290698
rect 371884 290634 371936 290640
rect 371700 290556 371752 290562
rect 371804 290550 371924 290578
rect 371700 290498 371752 290504
rect 371792 290488 371844 290494
rect 371792 290430 371844 290436
rect 371804 290193 371832 290430
rect 371790 290184 371846 290193
rect 371790 290119 371846 290128
rect 371700 289264 371752 289270
rect 371700 289206 371752 289212
rect 371712 289105 371740 289206
rect 371698 289096 371754 289105
rect 371698 289031 371754 289040
rect 371700 288584 371752 288590
rect 371698 288552 371700 288561
rect 371752 288552 371754 288561
rect 371698 288487 371754 288496
rect 371896 288153 371924 290550
rect 371882 288144 371938 288153
rect 371882 288079 371938 288088
rect 371988 286521 372016 414582
rect 372066 412584 372122 412593
rect 372066 412519 372068 412528
rect 372120 412519 372122 412528
rect 372068 412490 372120 412496
rect 372250 298072 372306 298081
rect 372250 298007 372306 298016
rect 372160 295996 372212 296002
rect 372160 295938 372212 295944
rect 372066 295352 372122 295361
rect 372066 295287 372122 295296
rect 372080 287054 372108 295287
rect 372172 295089 372200 295938
rect 372158 295080 372214 295089
rect 372158 295015 372214 295024
rect 372264 291786 372292 298007
rect 372342 296168 372398 296177
rect 372342 296103 372344 296112
rect 372396 296103 372398 296112
rect 372344 296074 372396 296080
rect 372540 291938 372568 429150
rect 372620 425060 372672 425066
rect 372620 425002 372672 425008
rect 372632 424425 372660 425002
rect 372618 424416 372674 424425
rect 372618 424351 372674 424360
rect 372632 369714 372660 424351
rect 372816 413137 372844 486934
rect 372908 485314 372936 556242
rect 373000 511222 373028 567870
rect 373264 565888 373316 565894
rect 373264 565830 373316 565836
rect 373276 556102 373304 565830
rect 373264 556096 373316 556102
rect 373264 556038 373316 556044
rect 372988 511216 373040 511222
rect 372988 511158 373040 511164
rect 372896 485308 372948 485314
rect 372896 485250 372948 485256
rect 372802 413128 372858 413137
rect 372802 413063 372858 413072
rect 372816 412634 372844 413063
rect 372724 412606 372844 412634
rect 372620 369708 372672 369714
rect 372620 369650 372672 369656
rect 372620 369572 372672 369578
rect 372620 369514 372672 369520
rect 372632 369170 372660 369514
rect 372620 369164 372672 369170
rect 372620 369106 372672 369112
rect 372620 350940 372672 350946
rect 372620 350882 372672 350888
rect 372356 291910 372568 291938
rect 372252 291780 372304 291786
rect 372252 291722 372304 291728
rect 372080 287026 372292 287054
rect 371974 286512 372030 286521
rect 371974 286447 372030 286456
rect 371608 286408 371660 286414
rect 371608 286350 371660 286356
rect 371516 286340 371568 286346
rect 371516 286282 371568 286288
rect 371146 285968 371202 285977
rect 371146 285903 371202 285912
rect 371056 247716 371108 247722
rect 371056 247658 371108 247664
rect 371068 247110 371096 247658
rect 370504 247104 370556 247110
rect 370504 247046 370556 247052
rect 371056 247104 371108 247110
rect 371056 247046 371108 247052
rect 370516 224262 370544 247046
rect 371160 229770 371188 285903
rect 371988 285734 372016 286447
rect 371976 285728 372028 285734
rect 371976 285670 372028 285676
rect 372264 284374 372292 287026
rect 372356 285433 372384 291910
rect 372436 291780 372488 291786
rect 372436 291722 372488 291728
rect 372342 285424 372398 285433
rect 372342 285359 372398 285368
rect 372448 284889 372476 291722
rect 372434 284880 372490 284889
rect 372434 284815 372490 284824
rect 372252 284368 372304 284374
rect 372250 284336 372252 284345
rect 372304 284336 372306 284345
rect 372250 284271 372306 284280
rect 371516 283620 371568 283626
rect 371516 283562 371568 283568
rect 371528 283257 371556 283562
rect 371514 283248 371570 283257
rect 371514 283183 371570 283192
rect 371606 282704 371662 282713
rect 371606 282639 371662 282648
rect 371620 282266 371648 282639
rect 371700 282328 371752 282334
rect 371700 282270 371752 282276
rect 371608 282260 371660 282266
rect 371608 282202 371660 282208
rect 371516 282192 371568 282198
rect 371712 282169 371740 282270
rect 371516 282134 371568 282140
rect 371698 282160 371754 282169
rect 371528 281625 371556 282134
rect 371698 282095 371754 282104
rect 371238 281616 371294 281625
rect 371238 281551 371294 281560
rect 371514 281616 371570 281625
rect 371514 281551 371570 281560
rect 371148 229764 371200 229770
rect 371148 229706 371200 229712
rect 371160 225622 371188 229706
rect 371252 225729 371280 281551
rect 371514 281072 371570 281081
rect 371514 281007 371570 281016
rect 371528 280838 371556 281007
rect 371516 280832 371568 280838
rect 371516 280774 371568 280780
rect 371528 280106 371556 280774
rect 371344 280078 371556 280106
rect 371238 225720 371294 225729
rect 371238 225655 371294 225664
rect 371148 225616 371200 225622
rect 371148 225558 371200 225564
rect 371344 224330 371372 280078
rect 371422 279984 371478 279993
rect 371422 279919 371478 279928
rect 371436 279478 371464 279919
rect 371424 279472 371476 279478
rect 371424 279414 371476 279420
rect 371606 279440 371662 279449
rect 371606 279375 371608 279384
rect 371660 279375 371662 279384
rect 371608 279346 371660 279352
rect 371606 278352 371662 278361
rect 371606 278287 371608 278296
rect 371660 278287 371662 278296
rect 371608 278258 371660 278264
rect 371422 277400 371478 277409
rect 371422 277335 371478 277344
rect 371436 276214 371464 277335
rect 372434 276312 372490 276321
rect 372434 276247 372436 276256
rect 372488 276247 372490 276256
rect 372436 276218 372488 276224
rect 371424 276208 371476 276214
rect 371424 276150 371476 276156
rect 371608 275800 371660 275806
rect 371606 275768 371608 275777
rect 371660 275768 371662 275777
rect 371606 275703 371662 275712
rect 372160 275256 372212 275262
rect 372158 275224 372160 275233
rect 372212 275224 372214 275233
rect 372158 275159 372214 275168
rect 371514 274136 371570 274145
rect 371514 274071 371570 274080
rect 371528 273290 371556 274071
rect 371608 273624 371660 273630
rect 371606 273592 371608 273601
rect 371660 273592 371662 273601
rect 371606 273527 371662 273536
rect 372632 273290 372660 350882
rect 372724 342922 372752 412606
rect 372908 412554 372936 485250
rect 373000 425066 373028 511158
rect 373276 505510 373304 556038
rect 373264 505504 373316 505510
rect 373264 505446 373316 505452
rect 373080 504212 373132 504218
rect 373080 504154 373132 504160
rect 372988 425060 373040 425066
rect 372988 425002 373040 425008
rect 373092 421297 373120 504154
rect 373264 500336 373316 500342
rect 373264 500278 373316 500284
rect 373276 455462 373304 500278
rect 373264 455456 373316 455462
rect 373264 455398 373316 455404
rect 373908 455456 373960 455462
rect 373908 455398 373960 455404
rect 373078 421288 373134 421297
rect 373078 421223 373134 421232
rect 373920 419830 373948 455398
rect 374012 436830 374040 581062
rect 378232 581052 378284 581058
rect 378232 580994 378284 581000
rect 377036 579828 377088 579834
rect 377036 579770 377088 579776
rect 375472 578332 375524 578338
rect 375472 578274 375524 578280
rect 375380 571532 375432 571538
rect 375380 571474 375432 571480
rect 374644 567724 374696 567730
rect 374644 567666 374696 567672
rect 374184 566228 374236 566234
rect 374184 566170 374236 566176
rect 374092 558204 374144 558210
rect 374092 558146 374144 558152
rect 374104 490346 374132 558146
rect 374196 506530 374224 566170
rect 374276 564732 374328 564738
rect 374276 564674 374328 564680
rect 374184 506524 374236 506530
rect 374184 506466 374236 506472
rect 374288 503198 374316 564674
rect 374368 563100 374420 563106
rect 374368 563042 374420 563048
rect 374276 503192 374328 503198
rect 374276 503134 374328 503140
rect 374092 490340 374144 490346
rect 374092 490282 374144 490288
rect 374000 436824 374052 436830
rect 374000 436766 374052 436772
rect 374092 421592 374144 421598
rect 374092 421534 374144 421540
rect 373908 419824 373960 419830
rect 373908 419766 373960 419772
rect 373356 419484 373408 419490
rect 373356 419426 373408 419432
rect 373264 418124 373316 418130
rect 373264 418066 373316 418072
rect 372896 412548 372948 412554
rect 372896 412490 372948 412496
rect 372908 393314 372936 412490
rect 372816 393286 372936 393314
rect 372712 342916 372764 342922
rect 372712 342858 372764 342864
rect 372816 341737 372844 393286
rect 372896 369708 372948 369714
rect 372896 369650 372948 369656
rect 372908 367538 372936 369650
rect 372896 367532 372948 367538
rect 372896 367474 372948 367480
rect 373276 354482 373304 418066
rect 373368 359174 373396 419426
rect 374000 369300 374052 369306
rect 374000 369242 374052 369248
rect 374012 367198 374040 369242
rect 374000 367192 374052 367198
rect 374000 367134 374052 367140
rect 374000 364812 374052 364818
rect 374000 364754 374052 364760
rect 373356 359168 373408 359174
rect 373356 359110 373408 359116
rect 373356 357876 373408 357882
rect 373356 357818 373408 357824
rect 373264 354476 373316 354482
rect 373264 354418 373316 354424
rect 373080 345228 373132 345234
rect 373080 345170 373132 345176
rect 372802 341728 372858 341737
rect 372802 341663 372858 341672
rect 372816 277394 372844 341663
rect 372986 278080 373042 278089
rect 372986 278015 373042 278024
rect 372724 277366 372844 277394
rect 371516 273284 371568 273290
rect 371516 273226 371568 273232
rect 372620 273284 372672 273290
rect 372620 273226 372672 273232
rect 371698 273048 371754 273057
rect 371698 272983 371754 272992
rect 371712 271794 371740 272983
rect 371882 272504 371938 272513
rect 371882 272439 371938 272448
rect 371790 271960 371846 271969
rect 371790 271895 371846 271904
rect 371700 271788 371752 271794
rect 371700 271730 371752 271736
rect 371424 269816 371476 269822
rect 371424 269758 371476 269764
rect 371436 269249 371464 269758
rect 371422 269240 371478 269249
rect 371422 269175 371478 269184
rect 371332 224324 371384 224330
rect 371332 224266 371384 224272
rect 370504 224256 370556 224262
rect 370504 224198 370556 224204
rect 370962 217424 371018 217433
rect 370962 217359 370964 217368
rect 371016 217359 371018 217368
rect 370964 217330 371016 217336
rect 370964 216232 371016 216238
rect 370962 216200 370964 216209
rect 371016 216200 371018 216209
rect 370962 216135 371018 216144
rect 370686 215112 370742 215121
rect 370686 215047 370688 215056
rect 370740 215047 370742 215056
rect 370688 215018 370740 215024
rect 370962 213888 371018 213897
rect 370962 213823 370964 213832
rect 371016 213823 371018 213832
rect 370964 213794 371016 213800
rect 370964 211608 371016 211614
rect 370962 211576 370964 211585
rect 371016 211576 371018 211585
rect 370962 211511 371018 211520
rect 370962 210488 371018 210497
rect 370962 210423 371018 210432
rect 370976 210322 371004 210423
rect 370964 210316 371016 210322
rect 370964 210258 371016 210264
rect 370962 209264 371018 209273
rect 370962 209199 370964 209208
rect 371016 209199 371018 209208
rect 370964 209170 371016 209176
rect 370962 208176 371018 208185
rect 370962 208111 370964 208120
rect 371016 208111 371018 208120
rect 370964 208082 371016 208088
rect 371238 205864 371294 205873
rect 371238 205799 371294 205808
rect 370962 197704 371018 197713
rect 370962 197639 370964 197648
rect 371016 197639 371018 197648
rect 370964 197610 371016 197616
rect 371148 197260 371200 197266
rect 371148 197202 371200 197208
rect 370870 196616 370926 196625
rect 370870 196551 370926 196560
rect 370504 156188 370556 156194
rect 370504 156130 370556 156136
rect 370410 149968 370466 149977
rect 370410 149903 370466 149912
rect 370318 148880 370374 148889
rect 370318 148815 370374 148824
rect 370226 141944 370282 141953
rect 370226 141879 370282 141888
rect 370516 140321 370544 156130
rect 370596 156120 370648 156126
rect 370596 156062 370648 156068
rect 370608 140865 370636 156062
rect 370594 140856 370650 140865
rect 370594 140791 370650 140800
rect 370502 140312 370558 140321
rect 370502 140247 370558 140256
rect 370134 139768 370190 139777
rect 370134 139703 370190 139712
rect 370042 133648 370098 133657
rect 370042 133583 370098 133592
rect 369858 132424 369914 132433
rect 369858 132359 369914 132368
rect 369490 132016 369546 132025
rect 369490 131951 369546 131960
rect 369398 131472 369454 131481
rect 369398 131407 369454 131416
rect 370044 130484 370096 130490
rect 370044 130426 370096 130432
rect 370056 130257 370084 130426
rect 370320 130416 370372 130422
rect 370320 130358 370372 130364
rect 370042 130248 370098 130257
rect 370042 130183 370098 130192
rect 369858 129160 369914 129169
rect 369858 129095 369914 129104
rect 369306 128616 369362 128625
rect 369306 128551 369362 128560
rect 369320 125458 369348 128551
rect 369398 126440 369454 126449
rect 369398 126375 369454 126384
rect 369308 125452 369360 125458
rect 369308 125394 369360 125400
rect 369320 125050 369348 125394
rect 369308 125044 369360 125050
rect 369308 124986 369360 124992
rect 360580 124766 360962 124794
rect 368966 124766 369164 124794
rect 362788 124086 362894 124114
rect 364918 124086 365208 124114
rect 362788 124001 362816 124086
rect 365180 124001 365208 124086
rect 362774 123992 362830 124001
rect 362774 123927 362830 123936
rect 365166 123992 365222 124001
rect 365166 123927 365222 123936
rect 366928 122126 366956 124100
rect 369412 124098 369440 126375
rect 369872 125186 369900 129095
rect 369950 128616 370006 128625
rect 369950 128551 370006 128560
rect 369964 125254 369992 128551
rect 369952 125248 370004 125254
rect 369952 125190 370004 125196
rect 369860 125180 369912 125186
rect 369860 125122 369912 125128
rect 370056 125118 370084 130183
rect 370332 130121 370360 130358
rect 370318 130112 370374 130121
rect 370318 130047 370374 130056
rect 370226 127936 370282 127945
rect 370226 127871 370282 127880
rect 370134 127392 370190 127401
rect 370134 127327 370190 127336
rect 370044 125112 370096 125118
rect 370044 125054 370096 125060
rect 369860 124772 369912 124778
rect 369860 124714 369912 124720
rect 369872 124409 369900 124714
rect 369858 124400 369914 124409
rect 369858 124335 369914 124344
rect 368204 124092 368256 124098
rect 368204 124034 368256 124040
rect 369400 124092 369452 124098
rect 369400 124034 369452 124040
rect 366916 122120 366968 122126
rect 366916 122062 366968 122068
rect 368216 117298 368244 124034
rect 369872 123486 369900 124335
rect 369950 123992 370006 124001
rect 369950 123927 370006 123936
rect 369860 123480 369912 123486
rect 369860 123422 369912 123428
rect 369964 122834 369992 123927
rect 369872 122806 369992 122834
rect 368204 117292 368256 117298
rect 368204 117234 368256 117240
rect 369872 102134 369900 122806
rect 370148 120086 370176 127327
rect 370240 124914 370268 127871
rect 370332 124982 370360 130047
rect 370410 126304 370466 126313
rect 370410 126239 370466 126248
rect 370424 125934 370452 126239
rect 370412 125928 370464 125934
rect 370412 125870 370464 125876
rect 370320 124976 370372 124982
rect 370320 124918 370372 124924
rect 370228 124908 370280 124914
rect 370228 124850 370280 124856
rect 370424 123554 370452 125870
rect 370502 125760 370558 125769
rect 370502 125695 370558 125704
rect 370412 123548 370464 123554
rect 370412 123490 370464 123496
rect 370136 120080 370188 120086
rect 370136 120022 370188 120028
rect 370516 111790 370544 125695
rect 370884 124914 370912 196551
rect 371056 193248 371108 193254
rect 371056 193190 371108 193196
rect 370964 191820 371016 191826
rect 370964 191762 371016 191768
rect 370976 156058 371004 191762
rect 371068 156194 371096 193190
rect 371056 156188 371108 156194
rect 371056 156130 371108 156136
rect 371160 156126 371188 197202
rect 371252 170542 371280 205799
rect 371330 202328 371386 202337
rect 371330 202263 371386 202272
rect 371240 170536 371292 170542
rect 371240 170478 371292 170484
rect 371240 170400 371292 170406
rect 371240 170342 371292 170348
rect 371252 164218 371280 170342
rect 371240 164212 371292 164218
rect 371240 164154 371292 164160
rect 371148 156120 371200 156126
rect 371148 156062 371200 156068
rect 370964 156052 371016 156058
rect 370964 155994 371016 156000
rect 371240 153060 371292 153066
rect 371240 153002 371292 153008
rect 371252 152969 371280 153002
rect 371238 152960 371294 152969
rect 371238 152895 371294 152904
rect 371240 152720 371292 152726
rect 371240 152662 371292 152668
rect 371252 149433 371280 152662
rect 371238 149424 371294 149433
rect 371238 149359 371294 149368
rect 371344 148458 371372 202263
rect 371436 198937 371464 269175
rect 371712 227714 371740 271730
rect 371804 271726 371832 271895
rect 371896 271862 371924 272439
rect 371884 271856 371936 271862
rect 371884 271798 371936 271804
rect 372252 271856 372304 271862
rect 372252 271798 372304 271804
rect 371792 271720 371844 271726
rect 371792 271662 371844 271668
rect 372160 271720 372212 271726
rect 372160 271662 372212 271668
rect 371790 270872 371846 270881
rect 371790 270807 371846 270816
rect 371804 270502 371832 270807
rect 371792 270496 371844 270502
rect 371792 270438 371844 270444
rect 372068 270496 372120 270502
rect 372068 270438 372120 270444
rect 371974 270328 372030 270337
rect 371974 270263 372030 270272
rect 371882 269784 371938 269793
rect 371882 269719 371938 269728
rect 371896 269074 371924 269719
rect 371884 269068 371936 269074
rect 371884 269010 371936 269016
rect 371712 227686 371832 227714
rect 371514 222048 371570 222057
rect 371514 221983 371570 221992
rect 371528 220794 371556 221983
rect 371516 220788 371568 220794
rect 371516 220730 371568 220736
rect 371804 206961 371832 227686
rect 371790 206952 371846 206961
rect 371790 206887 371846 206896
rect 371608 202360 371660 202366
rect 371608 202302 371660 202308
rect 371514 201240 371570 201249
rect 371514 201175 371570 201184
rect 371422 198928 371478 198937
rect 371422 198863 371478 198872
rect 371252 148430 371372 148458
rect 371252 126449 371280 148430
rect 371332 148300 371384 148306
rect 371332 148242 371384 148248
rect 371344 147801 371372 148242
rect 371330 147792 371386 147801
rect 371330 147727 371386 147736
rect 371332 147280 371384 147286
rect 371330 147248 371332 147257
rect 371384 147248 371386 147257
rect 371330 147183 371386 147192
rect 371332 145648 371384 145654
rect 371330 145616 371332 145625
rect 371384 145616 371386 145625
rect 371330 145551 371386 145560
rect 371332 145512 371384 145518
rect 371332 145454 371384 145460
rect 371344 145081 371372 145454
rect 371330 145072 371386 145081
rect 371330 145007 371386 145016
rect 371332 144560 371384 144566
rect 371330 144528 371332 144537
rect 371384 144528 371386 144537
rect 371330 144463 371386 144472
rect 371332 144152 371384 144158
rect 371330 144120 371332 144129
rect 371384 144120 371386 144129
rect 371330 144055 371386 144064
rect 371332 143472 371384 143478
rect 371332 143414 371384 143420
rect 371344 142497 371372 143414
rect 371330 142488 371386 142497
rect 371330 142423 371386 142432
rect 371332 139324 371384 139330
rect 371332 139266 371384 139272
rect 371344 138145 371372 139266
rect 371330 138136 371386 138145
rect 371330 138071 371386 138080
rect 371332 137624 371384 137630
rect 371330 137592 371332 137601
rect 371384 137592 371386 137601
rect 371330 137527 371386 137536
rect 371332 137352 371384 137358
rect 371332 137294 371384 137300
rect 371238 126440 371294 126449
rect 371238 126375 371294 126384
rect 371344 125934 371372 137294
rect 371332 125928 371384 125934
rect 371332 125870 371384 125876
rect 371436 125526 371464 198863
rect 371528 137358 371556 201175
rect 371620 200025 371648 202302
rect 371606 200016 371662 200025
rect 371606 199951 371662 199960
rect 371516 137352 371568 137358
rect 371516 137294 371568 137300
rect 371516 133000 371568 133006
rect 371516 132942 371568 132948
rect 371528 132841 371556 132942
rect 371514 132832 371570 132841
rect 371514 132767 371570 132776
rect 371620 126070 371648 199951
rect 371700 191820 371752 191826
rect 371700 191762 371752 191768
rect 371712 191146 371740 191762
rect 371700 191140 371752 191146
rect 371700 191082 371752 191088
rect 371700 169312 371752 169318
rect 371700 169254 371752 169260
rect 371712 169046 371740 169254
rect 371700 169040 371752 169046
rect 371700 168982 371752 168988
rect 371712 139398 371740 168982
rect 371700 139392 371752 139398
rect 371700 139334 371752 139340
rect 371700 139256 371752 139262
rect 371700 139198 371752 139204
rect 371712 138689 371740 139198
rect 371698 138680 371754 138689
rect 371698 138615 371754 138624
rect 371700 134360 371752 134366
rect 371698 134328 371700 134337
rect 371752 134328 371754 134337
rect 371698 134263 371754 134272
rect 371804 129033 371832 206887
rect 371896 202366 371924 269010
rect 371988 269006 372016 270263
rect 371976 269000 372028 269006
rect 371976 268942 372028 268948
rect 371884 202360 371936 202366
rect 371884 202302 371936 202308
rect 371988 201249 372016 268942
rect 372080 202337 372108 270438
rect 372172 204626 372200 271662
rect 372264 205873 372292 271798
rect 372526 271416 372582 271425
rect 372526 271351 372582 271360
rect 372540 270638 372568 271351
rect 372724 271266 372752 277366
rect 372804 275392 372856 275398
rect 372804 275334 372856 275340
rect 372816 274689 372844 275334
rect 372802 274680 372858 274689
rect 372802 274615 372858 274624
rect 372632 271238 372752 271266
rect 372528 270632 372580 270638
rect 372528 270574 372580 270580
rect 372540 269929 372568 270574
rect 372526 269920 372582 269929
rect 372526 269855 372582 269864
rect 372526 268696 372582 268705
rect 372632 268682 372660 271238
rect 372582 268654 372660 268682
rect 372526 268631 372582 268640
rect 372526 223136 372582 223145
rect 372526 223071 372582 223080
rect 372342 220824 372398 220833
rect 372342 220759 372398 220768
rect 372436 220788 372488 220794
rect 372250 205864 372306 205873
rect 372250 205799 372306 205808
rect 372250 204640 372306 204649
rect 372172 204598 372250 204626
rect 372250 204575 372306 204584
rect 372158 203552 372214 203561
rect 372158 203487 372214 203496
rect 372066 202328 372122 202337
rect 372066 202263 372122 202272
rect 371974 201240 372030 201249
rect 371974 201175 372030 201184
rect 371976 194472 372028 194478
rect 371976 194414 372028 194420
rect 371988 193254 372016 194414
rect 371976 193248 372028 193254
rect 371976 193190 372028 193196
rect 371884 170536 371936 170542
rect 371884 170478 371936 170484
rect 371896 167686 371924 170478
rect 371884 167680 371936 167686
rect 371884 167622 371936 167628
rect 371790 129024 371846 129033
rect 371790 128959 371846 128968
rect 371896 128625 371924 167622
rect 371976 166320 372028 166326
rect 371976 166262 372028 166268
rect 371988 163538 372016 166262
rect 371976 163532 372028 163538
rect 371976 163474 372028 163480
rect 372172 158817 372200 203487
rect 372264 161498 372292 204575
rect 372356 166326 372384 220759
rect 372436 220730 372488 220736
rect 372448 172582 372476 220730
rect 372436 172576 372488 172582
rect 372436 172518 372488 172524
rect 372448 169318 372476 172518
rect 372436 169312 372488 169318
rect 372436 169254 372488 169260
rect 372434 169008 372490 169017
rect 372540 168994 372568 223071
rect 372632 197674 372660 268654
rect 372816 258074 372844 274615
rect 372896 273284 372948 273290
rect 372896 273226 372948 273232
rect 372724 258046 372844 258074
rect 372724 210322 372752 258046
rect 372804 213920 372856 213926
rect 372804 213862 372856 213868
rect 372816 212809 372844 213862
rect 372802 212800 372858 212809
rect 372802 212735 372858 212744
rect 372712 210316 372764 210322
rect 372712 210258 372764 210264
rect 372620 197668 372672 197674
rect 372620 197610 372672 197616
rect 372816 176662 372844 212735
rect 372908 209234 372936 273226
rect 373000 217394 373028 278015
rect 373092 269006 373120 345170
rect 373276 313954 373304 354418
rect 373368 318918 373396 357818
rect 373356 318912 373408 318918
rect 373356 318854 373408 318860
rect 373816 318912 373868 318918
rect 373816 318854 373868 318860
rect 373264 313948 373316 313954
rect 373264 313890 373316 313896
rect 373276 275398 373304 313890
rect 373828 287054 373856 318854
rect 373828 287026 373948 287054
rect 373920 276282 373948 287026
rect 374012 279410 374040 364754
rect 374104 362506 374132 421534
rect 374288 420782 374316 503134
rect 374380 499662 374408 563042
rect 374460 562556 374512 562562
rect 374460 562498 374512 562504
rect 374368 499656 374420 499662
rect 374368 499598 374420 499604
rect 374276 420776 374328 420782
rect 374276 420718 374328 420724
rect 374184 419824 374236 419830
rect 374184 419766 374236 419772
rect 374092 362500 374144 362506
rect 374092 362442 374144 362448
rect 374000 279404 374052 279410
rect 374000 279346 374052 279352
rect 374104 278322 374132 362442
rect 374196 356794 374224 419766
rect 374288 419490 374316 420718
rect 374276 419484 374328 419490
rect 374276 419426 374328 419432
rect 374380 419234 374408 499598
rect 374472 498506 374500 562498
rect 374552 559156 374604 559162
rect 374552 559098 374604 559104
rect 374460 498500 374512 498506
rect 374460 498442 374512 498448
rect 374288 419206 374408 419234
rect 374288 419150 374316 419206
rect 374276 419144 374328 419150
rect 374276 419086 374328 419092
rect 374184 356788 374236 356794
rect 374184 356730 374236 356736
rect 374092 278316 374144 278322
rect 374092 278258 374144 278264
rect 373908 276276 373960 276282
rect 373908 276218 373960 276224
rect 373920 276026 373948 276218
rect 373920 275998 374132 276026
rect 373264 275392 373316 275398
rect 373264 275334 373316 275340
rect 373264 275256 373316 275262
rect 373264 275198 373316 275204
rect 373080 269000 373132 269006
rect 373080 268942 373132 268948
rect 372988 217388 373040 217394
rect 372988 217330 373040 217336
rect 373000 216714 373028 217330
rect 372988 216708 373040 216714
rect 372988 216650 373040 216656
rect 373276 213602 373304 275198
rect 373356 274644 373408 274650
rect 373356 274586 373408 274592
rect 373368 213926 373396 274586
rect 374000 273624 374052 273630
rect 374000 273566 374052 273572
rect 373540 216708 373592 216714
rect 373540 216650 373592 216656
rect 373356 213920 373408 213926
rect 373356 213862 373408 213868
rect 373276 213574 373488 213602
rect 373460 211614 373488 213574
rect 373448 211608 373500 211614
rect 373448 211550 373500 211556
rect 373264 210316 373316 210322
rect 373264 210258 373316 210264
rect 372896 209228 372948 209234
rect 372896 209170 372948 209176
rect 372908 208418 372936 209170
rect 372896 208412 372948 208418
rect 372896 208354 372948 208360
rect 372804 176656 372856 176662
rect 372804 176598 372856 176604
rect 372490 168966 372568 168994
rect 372434 168943 372490 168952
rect 372344 166320 372396 166326
rect 372344 166262 372396 166268
rect 372344 163532 372396 163538
rect 372344 163474 372396 163480
rect 372252 161492 372304 161498
rect 372252 161434 372304 161440
rect 372158 158808 372214 158817
rect 372158 158743 372214 158752
rect 371976 146872 372028 146878
rect 371976 146814 372028 146820
rect 371988 146713 372016 146814
rect 371974 146704 372030 146713
rect 371974 146639 372030 146648
rect 371976 146260 372028 146266
rect 371976 146202 372028 146208
rect 371988 146169 372016 146202
rect 371974 146160 372030 146169
rect 371974 146095 372030 146104
rect 371976 143064 372028 143070
rect 371974 143032 371976 143041
rect 372028 143032 372030 143041
rect 371974 142967 372030 142976
rect 372264 142154 372292 161434
rect 372080 142126 372292 142154
rect 371976 142112 372028 142118
rect 371976 142054 372028 142060
rect 371988 141409 372016 142054
rect 371974 141400 372030 141409
rect 371974 141335 372030 141344
rect 371976 139392 372028 139398
rect 371976 139334 372028 139340
rect 371988 135969 372016 139334
rect 371974 135960 372030 135969
rect 371974 135895 372030 135904
rect 371882 128616 371938 128625
rect 371882 128551 371938 128560
rect 372080 127945 372108 142126
rect 372160 139392 372212 139398
rect 372160 139334 372212 139340
rect 372172 139233 372200 139334
rect 372158 139224 372214 139233
rect 372158 139159 372214 139168
rect 372356 135425 372384 163474
rect 372448 153202 372476 168943
rect 373276 160750 373304 210258
rect 373356 208412 373408 208418
rect 373356 208354 373408 208360
rect 373368 165578 373396 208354
rect 373460 171834 373488 211550
rect 373552 178702 373580 216650
rect 374012 208146 374040 273566
rect 374104 229094 374132 275998
rect 374196 275806 374224 356730
rect 374288 355570 374316 419086
rect 374472 418198 374500 498442
rect 374564 492386 374592 559098
rect 374656 510066 374684 567666
rect 374644 510060 374696 510066
rect 374644 510002 374696 510008
rect 374920 510060 374972 510066
rect 374920 510002 374972 510008
rect 374828 506524 374880 506530
rect 374828 506466 374880 506472
rect 374552 492380 374604 492386
rect 374552 492322 374604 492328
rect 374552 490340 374604 490346
rect 374552 490282 374604 490288
rect 374460 418192 374512 418198
rect 374460 418134 374512 418140
rect 374564 414798 374592 490282
rect 374736 424720 374788 424726
rect 374736 424662 374788 424668
rect 374644 422612 374696 422618
rect 374644 422554 374696 422560
rect 374552 414792 374604 414798
rect 374552 414734 374604 414740
rect 374564 412634 374592 414734
rect 374472 412606 374592 412634
rect 374276 355564 374328 355570
rect 374276 355506 374328 355512
rect 374184 275800 374236 275806
rect 374184 275742 374236 275748
rect 374196 274650 374224 275742
rect 374288 275262 374316 355506
rect 374368 352164 374420 352170
rect 374368 352106 374420 352112
rect 374276 275256 374328 275262
rect 374276 275198 374328 275204
rect 374184 274644 374236 274650
rect 374184 274586 374236 274592
rect 374380 273630 374408 352106
rect 374472 346322 374500 412606
rect 374656 367810 374684 422554
rect 374748 369374 374776 424662
rect 374840 421598 374868 506466
rect 374932 423842 374960 510002
rect 375392 426426 375420 571474
rect 375484 434586 375512 578274
rect 376760 577040 376812 577046
rect 376760 576982 376812 576988
rect 376208 570308 376260 570314
rect 376208 570250 376260 570256
rect 376024 570036 376076 570042
rect 376024 569978 376076 569984
rect 375564 560924 375616 560930
rect 375564 560866 375616 560872
rect 375576 494834 375604 560866
rect 375656 558068 375708 558074
rect 375656 558010 375708 558016
rect 375564 494828 375616 494834
rect 375564 494770 375616 494776
rect 375564 494012 375616 494018
rect 375564 493954 375616 493960
rect 375472 434580 375524 434586
rect 375472 434522 375524 434528
rect 375380 426420 375432 426426
rect 375380 426362 375432 426368
rect 375472 426080 375524 426086
rect 375472 426022 375524 426028
rect 374920 423836 374972 423842
rect 374920 423778 374972 423784
rect 374828 421592 374880 421598
rect 374828 421534 374880 421540
rect 374736 369368 374788 369374
rect 374736 369310 374788 369316
rect 374644 367804 374696 367810
rect 374644 367746 374696 367752
rect 374932 366518 374960 423778
rect 375012 421660 375064 421666
rect 375012 421602 375064 421608
rect 374920 366512 374972 366518
rect 374920 366454 374972 366460
rect 375024 364818 375052 421602
rect 375288 369232 375340 369238
rect 375288 369174 375340 369180
rect 375300 368558 375328 369174
rect 375288 368552 375340 368558
rect 375288 368494 375340 368500
rect 375012 364812 375064 364818
rect 375012 364754 375064 364760
rect 374460 346316 374512 346322
rect 374460 346258 374512 346264
rect 374368 273624 374420 273630
rect 374368 273566 374420 273572
rect 374472 270502 374500 346258
rect 375288 299872 375340 299878
rect 375288 299814 375340 299820
rect 375196 298036 375248 298042
rect 375196 297978 375248 297984
rect 375208 297430 375236 297978
rect 375196 297424 375248 297430
rect 375196 297366 375248 297372
rect 375104 296744 375156 296750
rect 375104 296686 375156 296692
rect 375116 289921 375144 296686
rect 375102 289912 375158 289921
rect 375102 289847 375158 289856
rect 375208 289513 375236 297366
rect 375300 296206 375328 299814
rect 375288 296200 375340 296206
rect 375288 296142 375340 296148
rect 375194 289504 375250 289513
rect 375194 289439 375250 289448
rect 374552 285728 374604 285734
rect 374552 285670 374604 285676
rect 374460 270496 374512 270502
rect 374460 270438 374512 270444
rect 374564 240786 374592 285670
rect 375380 284368 375432 284374
rect 375380 284310 375432 284316
rect 374736 279404 374788 279410
rect 374736 279346 374788 279352
rect 374644 276208 374696 276214
rect 374644 276150 374696 276156
rect 374552 240780 374604 240786
rect 374552 240722 374604 240728
rect 374104 229066 374316 229094
rect 374184 218476 374236 218482
rect 374184 218418 374236 218424
rect 374000 208140 374052 208146
rect 374000 208082 374052 208088
rect 373632 179444 373684 179450
rect 373632 179386 373684 179392
rect 373540 178696 373592 178702
rect 373540 178638 373592 178644
rect 373448 171828 373500 171834
rect 373448 171770 373500 171776
rect 373356 165572 373408 165578
rect 373356 165514 373408 165520
rect 373264 160744 373316 160750
rect 373264 160686 373316 160692
rect 372620 153876 372672 153882
rect 372620 153818 372672 153824
rect 372632 153270 372660 153818
rect 372620 153264 372672 153270
rect 372620 153206 372672 153212
rect 372988 153264 373040 153270
rect 372988 153206 373040 153212
rect 372436 153196 372488 153202
rect 372436 153138 372488 153144
rect 372620 153128 372672 153134
rect 372620 153070 372672 153076
rect 372632 146962 372660 153070
rect 372712 152788 372764 152794
rect 372712 152730 372764 152736
rect 372724 152046 372752 152730
rect 372896 152516 372948 152522
rect 372896 152458 372948 152464
rect 372712 152040 372764 152046
rect 372712 151982 372764 151988
rect 372724 151814 372752 151982
rect 372908 151910 372936 152458
rect 372896 151904 372948 151910
rect 372896 151846 372948 151852
rect 372724 151786 372844 151814
rect 372632 146934 372752 146962
rect 372620 146804 372672 146810
rect 372620 146746 372672 146752
rect 372632 140418 372660 146746
rect 372620 140412 372672 140418
rect 372620 140354 372672 140360
rect 372724 137442 372752 146934
rect 372632 137414 372752 137442
rect 372342 135416 372398 135425
rect 372342 135351 372398 135360
rect 372526 133920 372582 133929
rect 372632 133906 372660 137414
rect 372816 137057 372844 151786
rect 372908 139398 372936 151846
rect 373000 143070 373028 153206
rect 372988 143064 373040 143070
rect 372988 143006 373040 143012
rect 372988 140412 373040 140418
rect 372988 140354 373040 140360
rect 372896 139392 372948 139398
rect 372896 139334 372948 139340
rect 372802 137048 372858 137057
rect 372802 136983 372858 136992
rect 372582 133878 372660 133906
rect 372526 133855 372582 133864
rect 373000 133006 373028 140354
rect 372988 133000 373040 133006
rect 372988 132942 373040 132948
rect 373276 130490 373304 160686
rect 373264 130484 373316 130490
rect 373264 130426 373316 130432
rect 373368 130422 373396 165514
rect 373460 151774 373488 171770
rect 373552 153134 373580 178638
rect 373644 154562 373672 179386
rect 373724 168360 373776 168366
rect 373724 168302 373776 168308
rect 373632 154556 373684 154562
rect 373632 154498 373684 154504
rect 373540 153128 373592 153134
rect 373540 153070 373592 153076
rect 373448 151768 373500 151774
rect 373448 151710 373500 151716
rect 373644 137630 373672 154498
rect 373736 153202 373764 168302
rect 373724 153196 373776 153202
rect 373724 153138 373776 153144
rect 373736 146810 373764 153138
rect 373724 146804 373776 146810
rect 373724 146746 373776 146752
rect 373632 137624 373684 137630
rect 373632 137566 373684 137572
rect 373356 130416 373408 130422
rect 373356 130358 373408 130364
rect 374012 129577 374040 208082
rect 374092 197668 374144 197674
rect 374092 197610 374144 197616
rect 373998 129568 374054 129577
rect 373998 129503 374054 129512
rect 372066 127936 372122 127945
rect 372066 127871 372122 127880
rect 371698 126440 371754 126449
rect 371698 126375 371754 126384
rect 371608 126064 371660 126070
rect 371608 126006 371660 126012
rect 371620 125769 371648 126006
rect 371712 126002 371740 126375
rect 371700 125996 371752 126002
rect 371700 125938 371752 125944
rect 371606 125760 371662 125769
rect 371606 125695 371662 125704
rect 371424 125520 371476 125526
rect 371424 125462 371476 125468
rect 371436 125225 371464 125462
rect 371422 125216 371478 125225
rect 371422 125151 371478 125160
rect 370872 124908 370924 124914
rect 370872 124850 370924 124856
rect 370884 124273 370912 124850
rect 370870 124264 370926 124273
rect 370870 124199 370926 124208
rect 370504 111784 370556 111790
rect 370504 111726 370556 111732
rect 371436 109002 371464 125151
rect 374104 124778 374132 197610
rect 374196 158710 374224 218418
rect 374288 213858 374316 229066
rect 374656 216238 374684 276150
rect 374748 220833 374776 279346
rect 374828 278316 374880 278322
rect 374828 278258 374880 278264
rect 374734 220824 374790 220833
rect 374734 220759 374790 220768
rect 374840 218482 374868 278258
rect 375102 231840 375158 231849
rect 375102 231775 375158 231784
rect 375116 226234 375144 231775
rect 375194 231704 375250 231713
rect 375194 231639 375250 231648
rect 375208 226302 375236 231639
rect 375196 226296 375248 226302
rect 375196 226238 375248 226244
rect 375104 226228 375156 226234
rect 375104 226170 375156 226176
rect 374828 218476 374880 218482
rect 374828 218418 374880 218424
rect 374644 216232 374696 216238
rect 374644 216174 374696 216180
rect 374368 215076 374420 215082
rect 374368 215018 374420 215024
rect 374276 213852 374328 213858
rect 374276 213794 374328 213800
rect 374184 158704 374236 158710
rect 374184 158646 374236 158652
rect 374196 158030 374224 158646
rect 374184 158024 374236 158030
rect 374184 157966 374236 157972
rect 374196 134366 374224 157966
rect 374288 156670 374316 213794
rect 374380 168366 374408 215018
rect 374460 189780 374512 189786
rect 374460 189722 374512 189728
rect 374368 168360 374420 168366
rect 374368 168302 374420 168308
rect 374276 156664 374328 156670
rect 374276 156606 374328 156612
rect 374472 144158 374500 189722
rect 374656 155242 374684 216174
rect 375392 194478 375420 284310
rect 375484 282334 375512 426022
rect 375576 416430 375604 493954
rect 375668 488102 375696 558010
rect 376036 556170 376064 569978
rect 376116 560380 376168 560386
rect 376116 560322 376168 560328
rect 376024 556164 376076 556170
rect 376024 556106 376076 556112
rect 375656 488096 375708 488102
rect 375656 488038 375708 488044
rect 375840 426624 375892 426630
rect 375840 426566 375892 426572
rect 375564 416424 375616 416430
rect 375564 416366 375616 416372
rect 375576 349858 375604 416366
rect 375656 412140 375708 412146
rect 375656 412082 375708 412088
rect 375564 349852 375616 349858
rect 375564 349794 375616 349800
rect 375564 347200 375616 347206
rect 375564 347142 375616 347148
rect 375472 282328 375524 282334
rect 375472 282270 375524 282276
rect 375576 270638 375604 347142
rect 375668 344010 375696 412082
rect 375656 344004 375708 344010
rect 375656 343946 375708 343952
rect 375564 270632 375616 270638
rect 375564 270574 375616 270580
rect 375668 269074 375696 343946
rect 375852 282266 375880 426566
rect 376036 426086 376064 556106
rect 376128 556034 376156 560322
rect 376116 556028 376168 556034
rect 376116 555970 376168 555976
rect 376128 494018 376156 555970
rect 376220 522986 376248 570250
rect 376208 522980 376260 522986
rect 376208 522922 376260 522928
rect 376668 522980 376720 522986
rect 376668 522922 376720 522928
rect 376680 522306 376708 522922
rect 376668 522300 376720 522306
rect 376668 522242 376720 522248
rect 376208 494828 376260 494834
rect 376208 494770 376260 494776
rect 376116 494012 376168 494018
rect 376116 493954 376168 493960
rect 376220 447166 376248 494770
rect 376208 447160 376260 447166
rect 376208 447102 376260 447108
rect 376680 442338 376708 522242
rect 376116 442332 376168 442338
rect 376116 442274 376168 442280
rect 376668 442332 376720 442338
rect 376668 442274 376720 442280
rect 376128 441658 376156 442274
rect 376116 441652 376168 441658
rect 376116 441594 376168 441600
rect 376128 426630 376156 441594
rect 376772 434654 376800 576982
rect 376944 575544 376996 575550
rect 376944 575486 376996 575492
rect 376852 569968 376904 569974
rect 376852 569910 376904 569916
rect 376760 434648 376812 434654
rect 376760 434590 376812 434596
rect 376864 427106 376892 569910
rect 376956 432818 376984 575486
rect 377048 437374 377076 579770
rect 378140 577516 378192 577522
rect 378140 577458 378192 577464
rect 378152 576978 378180 577458
rect 378140 576972 378192 576978
rect 378140 576914 378192 576920
rect 377128 558952 377180 558958
rect 377128 558894 377180 558900
rect 377140 493338 377168 558894
rect 377128 493332 377180 493338
rect 377128 493274 377180 493280
rect 377036 437368 377088 437374
rect 377036 437310 377088 437316
rect 376944 432812 376996 432818
rect 376944 432754 376996 432760
rect 376852 427100 376904 427106
rect 376852 427042 376904 427048
rect 376116 426624 376168 426630
rect 376116 426566 376168 426572
rect 376024 426080 376076 426086
rect 376024 426022 376076 426028
rect 376024 415676 376076 415682
rect 376024 415618 376076 415624
rect 376036 348702 376064 415618
rect 376116 413976 376168 413982
rect 376116 413918 376168 413924
rect 376024 348696 376076 348702
rect 376024 348638 376076 348644
rect 376036 309126 376064 348638
rect 376128 347206 376156 413918
rect 376864 412634 376892 427042
rect 377140 415682 377168 493274
rect 377220 492380 377272 492386
rect 377220 492322 377272 492328
rect 377128 415676 377180 415682
rect 377128 415618 377180 415624
rect 377232 413982 377260 492322
rect 377312 447160 377364 447166
rect 377312 447102 377364 447108
rect 377324 417450 377352 447102
rect 377496 442332 377548 442338
rect 377496 442274 377548 442280
rect 377508 433294 377536 442274
rect 378048 437368 378100 437374
rect 378048 437310 378100 437316
rect 378060 436762 378088 437310
rect 378048 436756 378100 436762
rect 378048 436698 378100 436704
rect 377496 433288 377548 433294
rect 377496 433230 377548 433236
rect 377404 432812 377456 432818
rect 377404 432754 377456 432760
rect 377312 417444 377364 417450
rect 377312 417386 377364 417392
rect 377220 413976 377272 413982
rect 377220 413918 377272 413924
rect 376772 412606 376892 412634
rect 376668 359304 376720 359310
rect 376668 359246 376720 359252
rect 376116 347200 376168 347206
rect 376116 347142 376168 347148
rect 376024 309120 376076 309126
rect 376024 309062 376076 309068
rect 376036 306374 376064 309062
rect 376036 306346 376248 306374
rect 375932 299124 375984 299130
rect 375932 299066 375984 299072
rect 375944 298382 375972 299066
rect 375932 298376 375984 298382
rect 375932 298318 375984 298324
rect 375944 288590 375972 298318
rect 376024 289808 376076 289814
rect 376024 289750 376076 289756
rect 376036 289270 376064 289750
rect 376024 289264 376076 289270
rect 376024 289206 376076 289212
rect 375932 288584 375984 288590
rect 375932 288526 375984 288532
rect 375840 282260 375892 282266
rect 375840 282202 375892 282208
rect 375944 277394 375972 288526
rect 375760 277366 375972 277394
rect 375656 269068 375708 269074
rect 375656 269010 375708 269016
rect 375472 236020 375524 236026
rect 375472 235962 375524 235968
rect 375380 194472 375432 194478
rect 375380 194414 375432 194420
rect 375288 189780 375340 189786
rect 375288 189722 375340 189728
rect 375300 189106 375328 189722
rect 375288 189100 375340 189106
rect 375288 189042 375340 189048
rect 374644 155236 374696 155242
rect 374644 155178 374696 155184
rect 374656 152590 374684 155178
rect 374644 152584 374696 152590
rect 374644 152526 374696 152532
rect 375484 148306 375512 235962
rect 375564 233300 375616 233306
rect 375564 233242 375616 233248
rect 375472 148300 375524 148306
rect 375472 148242 375524 148248
rect 375576 147286 375604 233242
rect 375656 231124 375708 231130
rect 375656 231066 375708 231072
rect 375668 230518 375696 231066
rect 375656 230512 375708 230518
rect 375656 230454 375708 230460
rect 375564 147280 375616 147286
rect 375564 147222 375616 147228
rect 375668 146878 375696 230454
rect 375760 225010 375788 277366
rect 376036 229094 376064 289206
rect 376116 278724 376168 278730
rect 376116 278666 376168 278672
rect 375852 229066 376064 229094
rect 375852 225078 375880 229066
rect 375840 225072 375892 225078
rect 375840 225014 375892 225020
rect 375748 225004 375800 225010
rect 375748 224946 375800 224952
rect 375656 146872 375708 146878
rect 375656 146814 375708 146820
rect 375760 144566 375788 224946
rect 375852 145518 375880 225014
rect 375932 223984 375984 223990
rect 375932 223926 375984 223932
rect 375944 145654 375972 223926
rect 376024 220924 376076 220930
rect 376024 220866 376076 220872
rect 376036 170406 376064 220866
rect 376128 220794 376156 278666
rect 376220 271726 376248 306346
rect 376680 299130 376708 359246
rect 376668 299124 376720 299130
rect 376668 299066 376720 299072
rect 376772 283626 376800 412606
rect 377036 366512 377088 366518
rect 377036 366454 377088 366460
rect 376760 283620 376812 283626
rect 376760 283562 376812 283568
rect 376944 283620 376996 283626
rect 376944 283562 376996 283568
rect 376852 282260 376904 282266
rect 376852 282202 376904 282208
rect 376208 271720 376260 271726
rect 376208 271662 376260 271668
rect 376668 233912 376720 233918
rect 376668 233854 376720 233860
rect 376680 233306 376708 233854
rect 376668 233300 376720 233306
rect 376668 233242 376720 233248
rect 376116 220788 376168 220794
rect 376116 220730 376168 220736
rect 376864 184890 376892 282202
rect 376956 187678 376984 283562
rect 377048 279478 377076 366454
rect 377324 354674 377352 417386
rect 377416 385694 377444 432754
rect 378152 432682 378180 576914
rect 378244 438190 378272 580994
rect 378784 580304 378836 580310
rect 378784 580246 378836 580252
rect 378796 579766 378824 580246
rect 378784 579760 378836 579766
rect 378784 579702 378836 579708
rect 378232 438184 378284 438190
rect 378232 438126 378284 438132
rect 378244 437510 378272 438126
rect 378232 437504 378284 437510
rect 378232 437446 378284 437452
rect 378796 436014 378824 579702
rect 380164 579692 380216 579698
rect 380164 579634 380216 579640
rect 379152 578264 379204 578270
rect 379152 578206 379204 578212
rect 379060 576904 379112 576910
rect 379060 576846 379112 576852
rect 378876 438932 378928 438938
rect 378876 438874 378928 438880
rect 378784 436008 378836 436014
rect 378784 435950 378836 435956
rect 378140 432676 378192 432682
rect 378140 432618 378192 432624
rect 378784 432676 378836 432682
rect 378784 432618 378836 432624
rect 377404 385688 377456 385694
rect 377404 385630 377456 385636
rect 377416 359310 377444 385630
rect 378796 371890 378824 432618
rect 378784 371884 378836 371890
rect 378784 371826 378836 371832
rect 377588 369368 377640 369374
rect 377588 369310 377640 369316
rect 377496 367804 377548 367810
rect 377496 367746 377548 367752
rect 377404 359304 377456 359310
rect 377404 359246 377456 359252
rect 377140 354646 377352 354674
rect 377140 351218 377168 354646
rect 377128 351212 377180 351218
rect 377128 351154 377180 351160
rect 377036 279472 377088 279478
rect 377036 279414 377088 279420
rect 377048 278730 377076 279414
rect 377036 278724 377088 278730
rect 377036 278666 377088 278672
rect 377140 271794 377168 351154
rect 377220 349852 377272 349858
rect 377220 349794 377272 349800
rect 377232 271862 377260 349794
rect 377312 342916 377364 342922
rect 377312 342858 377364 342864
rect 377220 271856 377272 271862
rect 377220 271798 377272 271804
rect 377128 271788 377180 271794
rect 377128 271730 377180 271736
rect 377324 270094 377352 342858
rect 377404 321632 377456 321638
rect 377404 321574 377456 321580
rect 377416 289814 377444 321574
rect 377404 289808 377456 289814
rect 377404 289750 377456 289756
rect 377404 286340 377456 286346
rect 377404 286282 377456 286288
rect 377312 270088 377364 270094
rect 377312 270030 377364 270036
rect 377416 242894 377444 286282
rect 377508 281518 377536 367746
rect 377600 282878 377628 369310
rect 378796 360262 378824 371826
rect 378048 360256 378100 360262
rect 378048 360198 378100 360204
rect 378784 360256 378836 360262
rect 378784 360198 378836 360204
rect 378060 322250 378088 360198
rect 378048 322244 378100 322250
rect 378048 322186 378100 322192
rect 378060 321638 378088 322186
rect 378048 321632 378100 321638
rect 378048 321574 378100 321580
rect 378784 314696 378836 314702
rect 378784 314638 378836 314644
rect 378232 291848 378284 291854
rect 378232 291790 378284 291796
rect 378140 289808 378192 289814
rect 378140 289750 378192 289756
rect 378152 289134 378180 289750
rect 378140 289128 378192 289134
rect 378140 289070 378192 289076
rect 377588 282872 377640 282878
rect 377588 282814 377640 282820
rect 378048 282872 378100 282878
rect 378048 282814 378100 282820
rect 377680 282328 377732 282334
rect 377680 282270 377732 282276
rect 377496 281512 377548 281518
rect 377496 281454 377548 281460
rect 377404 242888 377456 242894
rect 377404 242830 377456 242836
rect 376944 187672 376996 187678
rect 376944 187614 376996 187620
rect 376956 186998 376984 187614
rect 376944 186992 376996 186998
rect 376944 186934 376996 186940
rect 376852 184884 376904 184890
rect 376852 184826 376904 184832
rect 377692 182170 377720 282270
rect 378060 282198 378088 282814
rect 378048 282192 378100 282198
rect 378048 282134 378100 282140
rect 378048 281512 378100 281518
rect 378048 281454 378100 281460
rect 378060 280838 378088 281454
rect 378048 280832 378100 280838
rect 378048 280774 378100 280780
rect 377772 242888 377824 242894
rect 377772 242830 377824 242836
rect 377784 242214 377812 242830
rect 377772 242208 377824 242214
rect 377772 242150 377824 242156
rect 378152 224262 378180 289070
rect 378244 236706 378272 291790
rect 378796 289814 378824 314638
rect 378888 296546 378916 438874
rect 378968 437504 379020 437510
rect 378968 437446 379020 437452
rect 378876 296540 378928 296546
rect 378876 296482 378928 296488
rect 378888 295322 378916 296482
rect 378980 295390 379008 437446
rect 379072 434790 379100 576846
rect 379164 436150 379192 578206
rect 380176 437510 380204 579634
rect 380164 437504 380216 437510
rect 380164 437446 380216 437452
rect 379244 436824 379296 436830
rect 379244 436766 379296 436772
rect 379152 436144 379204 436150
rect 379152 436086 379204 436092
rect 379060 434784 379112 434790
rect 379060 434726 379112 434732
rect 379256 295458 379284 436766
rect 387064 436756 387116 436762
rect 387064 436698 387116 436704
rect 382924 436008 382976 436014
rect 382924 435950 382976 435956
rect 380164 434648 380216 434654
rect 380164 434590 380216 434596
rect 380176 384334 380204 434590
rect 381544 434580 381596 434586
rect 381544 434522 381596 434528
rect 380164 384328 380216 384334
rect 380164 384270 380216 384276
rect 380176 360262 380204 384270
rect 381556 369918 381584 434522
rect 382936 387122 382964 435950
rect 387076 398138 387104 436698
rect 395344 436144 395396 436150
rect 395344 436086 395396 436092
rect 393964 434784 394016 434790
rect 393964 434726 394016 434732
rect 387064 398132 387116 398138
rect 387064 398074 387116 398080
rect 382924 387116 382976 387122
rect 382924 387058 382976 387064
rect 383568 387116 383620 387122
rect 383568 387058 383620 387064
rect 381544 369912 381596 369918
rect 381544 369854 381596 369860
rect 382188 369912 382240 369918
rect 382188 369854 382240 369860
rect 379428 360256 379480 360262
rect 379428 360198 379480 360204
rect 380164 360256 380216 360262
rect 380164 360198 380216 360204
rect 379440 315314 379468 360198
rect 379428 315308 379480 315314
rect 379428 315250 379480 315256
rect 379440 314702 379468 315250
rect 379428 314696 379480 314702
rect 379428 314638 379480 314644
rect 379428 298784 379480 298790
rect 379428 298726 379480 298732
rect 379244 295452 379296 295458
rect 379244 295394 379296 295400
rect 378968 295384 379020 295390
rect 378968 295326 379020 295332
rect 378876 295316 378928 295322
rect 378876 295258 378928 295264
rect 378980 295254 379008 295326
rect 378968 295248 379020 295254
rect 378968 295190 379020 295196
rect 379256 293894 379284 295394
rect 379244 293888 379296 293894
rect 379244 293830 379296 293836
rect 379440 291854 379468 298726
rect 382200 298450 382228 369854
rect 382280 298852 382332 298858
rect 382280 298794 382332 298800
rect 382188 298444 382240 298450
rect 382188 298386 382240 298392
rect 379428 291848 379480 291854
rect 379428 291790 379480 291796
rect 382200 291174 382228 298386
rect 380900 291168 380952 291174
rect 380900 291110 380952 291116
rect 382188 291168 382240 291174
rect 382188 291110 382240 291116
rect 380912 290562 380940 291110
rect 380900 290556 380952 290562
rect 380900 290498 380952 290504
rect 378784 289808 378836 289814
rect 378784 289750 378836 289756
rect 378232 236700 378284 236706
rect 378232 236642 378284 236648
rect 378244 236026 378272 236642
rect 378232 236020 378284 236026
rect 378232 235962 378284 235968
rect 380912 231130 380940 290498
rect 382292 290494 382320 298794
rect 383580 298790 383608 387058
rect 387076 362982 387104 398074
rect 393976 394670 394004 434726
rect 395356 396030 395384 436086
rect 395344 396024 395396 396030
rect 395344 395966 395396 395972
rect 395988 396024 396040 396030
rect 395988 395966 396040 395972
rect 396000 395350 396028 395966
rect 395988 395344 396040 395350
rect 395988 395286 396040 395292
rect 393964 394664 394016 394670
rect 393964 394606 394016 394612
rect 394608 394664 394660 394670
rect 394608 394606 394660 394612
rect 394620 393990 394648 394606
rect 394608 393984 394660 393990
rect 394608 393926 394660 393932
rect 389088 367940 389140 367946
rect 389088 367882 389140 367888
rect 386328 362976 386380 362982
rect 386328 362918 386380 362924
rect 387064 362976 387116 362982
rect 387064 362918 387116 362924
rect 386340 310146 386368 362918
rect 385776 310140 385828 310146
rect 385776 310082 385828 310088
rect 386328 310140 386380 310146
rect 386328 310082 386380 310088
rect 383568 298784 383620 298790
rect 383568 298726 383620 298732
rect 385788 292534 385816 310082
rect 386340 309806 386368 310082
rect 386328 309800 386380 309806
rect 386328 309742 386380 309748
rect 389100 296682 389128 367882
rect 390468 367872 390520 367878
rect 390468 367814 390520 367820
rect 389088 296676 389140 296682
rect 389088 296618 389140 296624
rect 389100 296478 389128 296618
rect 390480 296614 390508 367814
rect 394620 298858 394648 393926
rect 396000 318782 396028 395286
rect 395344 318776 395396 318782
rect 395344 318718 395396 318724
rect 395988 318776 396040 318782
rect 395988 318718 396040 318724
rect 395356 318102 395384 318718
rect 395344 318096 395396 318102
rect 395344 318038 395396 318044
rect 394608 298852 394660 298858
rect 394608 298794 394660 298800
rect 390468 296608 390520 296614
rect 390468 296550 390520 296556
rect 389088 296472 389140 296478
rect 389088 296414 389140 296420
rect 390480 296138 390508 296550
rect 391940 296200 391992 296206
rect 391940 296142 391992 296148
rect 390468 296132 390520 296138
rect 390468 296074 390520 296080
rect 388444 296064 388496 296070
rect 388444 296006 388496 296012
rect 388456 295390 388484 296006
rect 388444 295384 388496 295390
rect 388444 295326 388496 295332
rect 385776 292528 385828 292534
rect 385776 292470 385828 292476
rect 386328 291848 386380 291854
rect 386328 291790 386380 291796
rect 386340 291242 386368 291790
rect 385684 291236 385736 291242
rect 385684 291178 385736 291184
rect 386328 291236 386380 291242
rect 386328 291178 386380 291184
rect 382280 290488 382332 290494
rect 382280 290430 382332 290436
rect 380900 231124 380952 231130
rect 380900 231066 380952 231072
rect 382292 227730 382320 290430
rect 385696 233918 385724 291178
rect 388456 249082 388484 295326
rect 388444 249076 388496 249082
rect 388444 249018 388496 249024
rect 385684 233912 385736 233918
rect 385684 233854 385736 233860
rect 382280 227724 382332 227730
rect 382280 227666 382332 227672
rect 382292 227050 382320 227666
rect 382280 227044 382332 227050
rect 382280 226986 382332 226992
rect 390480 224942 390508 296074
rect 391952 295866 391980 296142
rect 391940 295860 391992 295866
rect 391940 295802 391992 295808
rect 393228 295860 393280 295866
rect 393228 295802 393280 295808
rect 390468 224936 390520 224942
rect 390468 224878 390520 224884
rect 393240 224874 393268 295802
rect 395356 291854 395384 318038
rect 396736 307222 396764 699654
rect 425704 585268 425756 585274
rect 425704 585210 425756 585216
rect 425716 576162 425744 585210
rect 427820 583976 427872 583982
rect 427820 583918 427872 583924
rect 427832 580310 427860 583918
rect 427820 580304 427872 580310
rect 427820 580246 427872 580252
rect 425704 576156 425756 576162
rect 425704 576098 425756 576104
rect 399484 437504 399536 437510
rect 399484 437446 399536 437452
rect 399496 388482 399524 437446
rect 399484 388476 399536 388482
rect 399484 388418 399536 388424
rect 400128 388476 400180 388482
rect 400128 388418 400180 388424
rect 396724 307216 396776 307222
rect 396724 307158 396776 307164
rect 400140 298217 400168 388418
rect 429212 305794 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 699718 462360 703520
rect 478524 700534 478552 703520
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 461584 699712 461636 699718
rect 461584 699654 461636 699660
rect 462320 699712 462372 699718
rect 462320 699654 462372 699660
rect 445666 585440 445722 585449
rect 445722 585398 445800 585426
rect 445666 585375 445722 585384
rect 444746 584352 444802 584361
rect 444746 584287 444802 584296
rect 430580 584044 430632 584050
rect 430580 583986 430632 583992
rect 430592 577522 430620 583986
rect 444760 583914 444788 584287
rect 444748 583908 444800 583914
rect 444748 583850 444800 583856
rect 442998 583128 443054 583137
rect 442998 583063 443054 583072
rect 430580 577516 430632 577522
rect 430580 577458 430632 577464
rect 441618 577144 441674 577153
rect 441618 577079 441674 577088
rect 441632 576854 441660 577079
rect 441632 576826 441752 576854
rect 441618 559464 441674 559473
rect 441618 559399 441674 559408
rect 441632 558074 441660 559399
rect 441620 558068 441672 558074
rect 441620 558010 441672 558016
rect 441724 557534 441752 576826
rect 441802 573336 441858 573345
rect 441802 573271 441858 573280
rect 441632 557506 441752 557534
rect 441632 556102 441660 557506
rect 441710 556880 441766 556889
rect 441710 556815 441712 556824
rect 441764 556815 441766 556824
rect 441712 556786 441764 556792
rect 441620 556096 441672 556102
rect 431972 556022 432952 556050
rect 434884 556022 435220 556050
rect 431972 499574 432000 556022
rect 435192 554742 435220 556022
rect 436756 556022 436908 556050
rect 438932 556022 438992 556050
rect 440956 556022 441108 556050
rect 441620 556038 441672 556044
rect 435180 554736 435232 554742
rect 435180 554678 435232 554684
rect 435192 553489 435220 554678
rect 436756 553489 436784 556022
rect 438964 554062 438992 556022
rect 438952 554056 439004 554062
rect 438952 553998 439004 554004
rect 435178 553480 435234 553489
rect 435178 553415 435234 553424
rect 436742 553480 436798 553489
rect 436742 553415 436798 553424
rect 431972 499546 432552 499574
rect 432524 484106 432552 499546
rect 441080 484106 441108 556022
rect 441710 507376 441766 507385
rect 441710 507311 441766 507320
rect 441618 504656 441674 504665
rect 441618 504591 441674 504600
rect 432524 484078 433012 484106
rect 434884 484078 435220 484106
rect 432984 482798 433012 484078
rect 435192 483993 435220 484078
rect 436756 484078 436908 484106
rect 438932 484078 438992 484106
rect 440956 484078 441108 484106
rect 436756 483993 436784 484078
rect 435178 483984 435234 483993
rect 435178 483919 435234 483928
rect 436742 483984 436798 483993
rect 436742 483919 436798 483928
rect 435192 483002 435220 483919
rect 435180 482996 435232 483002
rect 435180 482938 435232 482944
rect 436756 482934 436784 483919
rect 436744 482928 436796 482934
rect 436744 482870 436796 482876
rect 432972 482792 433024 482798
rect 432972 482734 433024 482740
rect 438964 482390 438992 484078
rect 440988 482866 441016 484078
rect 440976 482860 441028 482866
rect 440976 482802 441028 482808
rect 438952 482384 439004 482390
rect 438952 482326 439004 482332
rect 432892 411998 432952 412026
rect 434884 411998 434944 412026
rect 432892 409766 432920 411998
rect 432880 409760 432932 409766
rect 432880 409702 432932 409708
rect 432892 408542 432920 409702
rect 434916 408649 434944 411998
rect 436848 411998 436908 412026
rect 438872 411998 438932 412026
rect 440956 411998 441108 412026
rect 436848 409834 436876 411998
rect 436836 409828 436888 409834
rect 436836 409770 436888 409776
rect 436848 408649 436876 409770
rect 438872 409154 438900 411998
rect 441080 409698 441108 411998
rect 441068 409692 441120 409698
rect 441068 409634 441120 409640
rect 441080 409601 441108 409634
rect 441066 409592 441122 409601
rect 441066 409527 441122 409536
rect 438860 409148 438912 409154
rect 438860 409090 438912 409096
rect 434902 408640 434958 408649
rect 434902 408575 434958 408584
rect 436834 408640 436890 408649
rect 436834 408575 436890 408584
rect 431960 408536 432012 408542
rect 431960 408478 432012 408484
rect 432880 408536 432932 408542
rect 432880 408478 432932 408484
rect 431972 364334 432000 408478
rect 441632 371890 441660 504591
rect 441724 387122 441752 507311
rect 441816 492561 441844 573271
rect 441894 567624 441950 567633
rect 441894 567559 441950 567568
rect 441802 492552 441858 492561
rect 441802 492487 441858 492496
rect 441908 489705 441936 567559
rect 441986 561776 442042 561785
rect 441986 561711 442042 561720
rect 441894 489696 441950 489705
rect 441894 489631 441950 489640
rect 441908 488578 441936 489631
rect 441896 488572 441948 488578
rect 441896 488514 441948 488520
rect 442000 486985 442028 561711
rect 442078 558920 442134 558929
rect 442078 558855 442134 558864
rect 441986 486976 442042 486985
rect 441986 486911 442042 486920
rect 442092 485217 442120 558855
rect 443012 496505 443040 583063
rect 443090 580816 443146 580825
rect 443090 580751 443146 580760
rect 442998 496496 443054 496505
rect 442998 496431 443054 496440
rect 443104 495417 443132 580751
rect 444746 579728 444802 579737
rect 444746 579663 444748 579672
rect 444800 579663 444802 579672
rect 444748 579634 444800 579640
rect 444930 578504 444986 578513
rect 444930 578439 444932 578448
rect 444984 578439 444986 578448
rect 444932 578410 444984 578416
rect 444746 576192 444802 576201
rect 444746 576127 444802 576136
rect 444760 575550 444788 576127
rect 444748 575544 444800 575550
rect 444748 575486 444800 575492
rect 444562 575104 444618 575113
rect 444562 575039 444618 575048
rect 444576 574122 444604 575039
rect 444564 574116 444616 574122
rect 444564 574058 444616 574064
rect 444838 571568 444894 571577
rect 444838 571503 444840 571512
rect 444892 571503 444894 571512
rect 444840 571474 444892 571480
rect 443182 570480 443238 570489
rect 443182 570415 443238 570424
rect 443090 495408 443146 495417
rect 443090 495343 443146 495352
rect 442906 494864 442962 494873
rect 442906 494799 442962 494808
rect 442920 494086 442948 494799
rect 442448 494080 442500 494086
rect 442448 494022 442500 494028
rect 442908 494080 442960 494086
rect 442908 494022 442960 494028
rect 442356 488572 442408 488578
rect 442356 488514 442408 488520
rect 442078 485208 442134 485217
rect 442078 485143 442134 485152
rect 442080 455456 442132 455462
rect 442080 455398 442132 455404
rect 441802 435568 441858 435577
rect 441802 435503 441858 435512
rect 441712 387116 441764 387122
rect 441712 387058 441764 387064
rect 441620 371884 441672 371890
rect 441620 371826 441672 371832
rect 441632 369594 441660 371826
rect 441540 369566 441660 369594
rect 441344 369232 441396 369238
rect 441344 369174 441396 369180
rect 441356 368937 441384 369174
rect 441342 368928 441398 368937
rect 441342 368863 441398 368872
rect 441540 368778 441568 369566
rect 441618 369472 441674 369481
rect 441618 369407 441674 369416
rect 441632 369306 441660 369407
rect 441620 369300 441672 369306
rect 441620 369242 441672 369248
rect 441540 368750 441660 368778
rect 441632 368098 441660 368750
rect 441540 368070 441660 368098
rect 441344 367872 441396 367878
rect 441342 367840 441344 367849
rect 441396 367840 441398 367849
rect 441342 367775 441398 367784
rect 441540 367690 441568 368070
rect 441620 367940 441672 367946
rect 441620 367882 441672 367888
rect 441632 367849 441660 367882
rect 441618 367840 441674 367849
rect 441618 367775 441674 367784
rect 441540 367662 441660 367690
rect 431972 364306 432552 364334
rect 432524 340082 432552 364306
rect 441632 361321 441660 367662
rect 441724 364041 441752 387058
rect 441710 364032 441766 364041
rect 441710 363967 441766 363976
rect 441618 361312 441674 361321
rect 441618 361247 441674 361256
rect 441816 354674 441844 435503
rect 441894 429312 441950 429321
rect 441894 429247 441950 429256
rect 441724 354646 441844 354674
rect 441724 351121 441752 354646
rect 441710 351112 441766 351121
rect 441710 351047 441766 351056
rect 441908 348537 441936 429247
rect 442092 428777 442120 455398
rect 442264 447160 442316 447166
rect 442264 447102 442316 447108
rect 442078 428768 442134 428777
rect 442078 428703 442134 428712
rect 441986 424008 442042 424017
rect 441986 423943 442042 423952
rect 441894 348528 441950 348537
rect 441894 348463 441950 348472
rect 441908 347750 441936 348463
rect 441896 347744 441948 347750
rect 441896 347686 441948 347692
rect 442000 345817 442028 423943
rect 442276 422929 442304 447102
rect 442368 424153 442396 488514
rect 442460 435713 442488 494022
rect 442998 493912 443054 493921
rect 442998 493847 443054 493856
rect 442538 492280 442594 492289
rect 442538 492215 442594 492224
rect 442446 435704 442502 435713
rect 442446 435639 442502 435648
rect 442552 429865 442580 492215
rect 442630 485752 442686 485761
rect 442630 485687 442686 485696
rect 442538 429856 442594 429865
rect 442538 429791 442594 429800
rect 442354 424144 442410 424153
rect 442354 424079 442410 424088
rect 442262 422920 442318 422929
rect 442262 422855 442318 422864
rect 442078 419520 442134 419529
rect 442078 419455 442134 419464
rect 441986 345808 442042 345817
rect 441986 345743 442042 345752
rect 441894 343632 441950 343641
rect 441894 343567 441950 343576
rect 441802 343088 441858 343097
rect 441802 343023 441858 343032
rect 441632 340950 441660 340981
rect 441620 340944 441672 340950
rect 441618 340912 441620 340921
rect 441672 340912 441674 340921
rect 441618 340847 441674 340856
rect 436558 340096 436614 340105
rect 432524 340054 432952 340082
rect 431866 338056 431922 338065
rect 431866 337991 431922 338000
rect 431774 337920 431830 337929
rect 431774 337855 431830 337864
rect 431224 337476 431276 337482
rect 431224 337418 431276 337424
rect 429200 305788 429252 305794
rect 429200 305730 429252 305736
rect 429844 298580 429896 298586
rect 429844 298522 429896 298528
rect 400126 298208 400182 298217
rect 400126 298143 400182 298152
rect 400140 293962 400168 298143
rect 425704 296812 425756 296818
rect 425704 296754 425756 296760
rect 400680 296132 400732 296138
rect 400680 296074 400732 296080
rect 400692 295458 400720 296074
rect 400680 295452 400732 295458
rect 400680 295394 400732 295400
rect 400128 293956 400180 293962
rect 400128 293898 400180 293904
rect 395344 291848 395396 291854
rect 395344 291790 395396 291796
rect 400692 287054 400720 295394
rect 400692 287026 400904 287054
rect 400876 246362 400904 287026
rect 425716 282878 425744 296754
rect 428464 295928 428516 295934
rect 428464 295870 428516 295876
rect 425704 282872 425756 282878
rect 425704 282814 425756 282820
rect 428476 281518 428504 295870
rect 428464 281512 428516 281518
rect 428464 281454 428516 281460
rect 429856 266218 429884 298522
rect 429844 266212 429896 266218
rect 429844 266154 429896 266160
rect 400864 246356 400916 246362
rect 400864 246298 400916 246304
rect 406384 240780 406436 240786
rect 406384 240722 406436 240728
rect 406396 240174 406424 240722
rect 406384 240168 406436 240174
rect 406384 240110 406436 240116
rect 394148 227044 394200 227050
rect 394148 226986 394200 226992
rect 394160 226370 394188 226986
rect 394148 226364 394200 226370
rect 394148 226306 394200 226312
rect 394608 226364 394660 226370
rect 394608 226306 394660 226312
rect 393228 224868 393280 224874
rect 393228 224810 393280 224816
rect 378140 224256 378192 224262
rect 378140 224198 378192 224204
rect 378152 223990 378180 224198
rect 378140 223984 378192 223990
rect 378140 223926 378192 223932
rect 381544 195356 381596 195362
rect 381544 195298 381596 195304
rect 378048 184884 378100 184890
rect 378048 184826 378100 184832
rect 378060 184210 378088 184826
rect 378048 184204 378100 184210
rect 378048 184146 378100 184152
rect 377680 182164 377732 182170
rect 377680 182106 377732 182112
rect 378048 182164 378100 182170
rect 378048 182106 378100 182112
rect 378060 181490 378088 182106
rect 378048 181484 378100 181490
rect 378048 181426 378100 181432
rect 376024 170400 376076 170406
rect 376024 170342 376076 170348
rect 375932 145648 375984 145654
rect 375932 145590 375984 145596
rect 375840 145512 375892 145518
rect 375840 145454 375892 145460
rect 375748 144560 375800 144566
rect 375748 144502 375800 144508
rect 374460 144152 374512 144158
rect 374460 144094 374512 144100
rect 381556 142118 381584 195298
rect 394620 156534 394648 226306
rect 399484 184204 399536 184210
rect 399484 184146 399536 184152
rect 395344 181484 395396 181490
rect 395344 181426 395396 181432
rect 393964 156528 394016 156534
rect 393964 156470 394016 156476
rect 394608 156528 394660 156534
rect 394608 156470 394660 156476
rect 393976 146266 394004 156470
rect 394620 156262 394648 156470
rect 394608 156256 394660 156262
rect 394608 156198 394660 156204
rect 393964 146260 394016 146266
rect 393964 146202 394016 146208
rect 381544 142112 381596 142118
rect 381544 142054 381596 142060
rect 395356 139330 395384 181426
rect 395344 139324 395396 139330
rect 395344 139266 395396 139272
rect 395988 139324 396040 139330
rect 395988 139266 396040 139272
rect 396000 138718 396028 139266
rect 399496 139262 399524 184146
rect 406396 143546 406424 240110
rect 406384 143540 406436 143546
rect 406384 143482 406436 143488
rect 399484 139256 399536 139262
rect 399484 139198 399536 139204
rect 399496 138786 399524 139198
rect 399484 138780 399536 138786
rect 399484 138722 399536 138728
rect 395988 138712 396040 138718
rect 395988 138654 396040 138660
rect 429844 138712 429896 138718
rect 429844 138654 429896 138660
rect 374184 134360 374236 134366
rect 374184 134302 374236 134308
rect 374828 125384 374880 125390
rect 374828 125326 374880 125332
rect 374840 124778 374868 125326
rect 429856 124778 429884 138654
rect 374092 124772 374144 124778
rect 374092 124714 374144 124720
rect 374828 124772 374880 124778
rect 374828 124714 374880 124720
rect 429844 124772 429896 124778
rect 429844 124714 429896 124720
rect 371424 108996 371476 109002
rect 371424 108938 371476 108944
rect 369860 102128 369912 102134
rect 369860 102070 369912 102076
rect 359464 99612 359516 99618
rect 359464 99554 359516 99560
rect 431236 99550 431264 337418
rect 431788 266354 431816 337855
rect 431776 266348 431828 266354
rect 431776 266290 431828 266296
rect 431880 266286 431908 337991
rect 432524 335354 432552 340054
rect 434870 339969 434898 340068
rect 440790 340096 440846 340105
rect 436614 340054 436908 340082
rect 438932 340054 438992 340082
rect 436558 340031 436614 340040
rect 434856 339960 434912 339969
rect 434856 339895 434912 339904
rect 434870 339810 434898 339895
rect 434824 339782 434898 339810
rect 434824 337929 434852 339782
rect 436572 338065 436600 340031
rect 436558 338056 436614 338065
rect 436558 337991 436614 338000
rect 434810 337920 434866 337929
rect 434810 337855 434866 337864
rect 438964 337482 438992 340054
rect 440846 340054 441108 340082
rect 440790 340031 440846 340040
rect 438952 337476 439004 337482
rect 438952 337418 439004 337424
rect 431972 335326 432552 335354
rect 431972 287054 432000 335326
rect 431972 287026 432552 287054
rect 432524 268546 432552 287026
rect 441080 268682 441108 340054
rect 441632 271561 441660 340847
rect 441710 296984 441766 296993
rect 441710 296919 441766 296928
rect 441724 296818 441752 296919
rect 441712 296812 441764 296818
rect 441712 296754 441764 296760
rect 441710 296032 441766 296041
rect 441710 295967 441766 295976
rect 441724 295934 441752 295967
rect 441712 295928 441764 295934
rect 441712 295870 441764 295876
rect 441816 275777 441844 343023
rect 441908 309126 441936 343567
rect 442092 343369 442120 419455
rect 442644 415993 442672 485687
rect 443012 433401 443040 493847
rect 443196 490657 443224 570415
rect 444930 569256 444986 569265
rect 444930 569191 444986 569200
rect 444944 568614 444972 569191
rect 444932 568608 444984 568614
rect 444932 568550 444984 568556
rect 443274 566944 443330 566953
rect 443274 566879 443330 566888
rect 443288 499574 443316 566879
rect 444470 565856 444526 565865
rect 444470 565791 444526 565800
rect 444378 564632 444434 564641
rect 444378 564567 444380 564576
rect 444432 564567 444434 564576
rect 444380 564538 444432 564544
rect 444378 561232 444434 561241
rect 444378 561167 444380 561176
rect 444432 561167 444434 561176
rect 444380 561138 444432 561144
rect 444378 557696 444434 557705
rect 444378 557631 444380 557640
rect 444432 557631 444434 557640
rect 444380 557602 444432 557608
rect 444484 556034 444512 565791
rect 445666 563544 445722 563553
rect 445666 563479 445722 563488
rect 445680 563106 445708 563479
rect 445668 563100 445720 563106
rect 445668 563042 445720 563048
rect 444472 556028 444524 556034
rect 444472 555970 444524 555976
rect 444380 513800 444432 513806
rect 444378 513768 444380 513777
rect 444932 513800 444984 513806
rect 444432 513768 444434 513777
rect 444932 513742 444984 513748
rect 444378 513703 444434 513712
rect 444838 513224 444894 513233
rect 444838 513159 444894 513168
rect 444564 512780 444616 512786
rect 444564 512722 444616 512728
rect 444378 512680 444434 512689
rect 444378 512615 444434 512624
rect 443288 499546 443500 499574
rect 443182 490648 443238 490657
rect 443182 490583 443238 490592
rect 443196 489914 443224 490583
rect 443104 489886 443224 489914
rect 443104 488782 443132 489886
rect 443472 489025 443500 499546
rect 443826 496496 443882 496505
rect 443826 496431 443882 496440
rect 443642 495408 443698 495417
rect 443642 495343 443698 495352
rect 443550 491736 443606 491745
rect 443550 491671 443606 491680
rect 443564 491366 443592 491671
rect 443552 491360 443604 491366
rect 443552 491302 443604 491308
rect 443458 489016 443514 489025
rect 443458 488951 443514 488960
rect 443092 488776 443144 488782
rect 443092 488718 443144 488724
rect 443274 486432 443330 486441
rect 443274 486367 443330 486376
rect 442998 433392 443054 433401
rect 442998 433327 443054 433336
rect 442170 415984 442226 415993
rect 442170 415919 442226 415928
rect 442630 415984 442686 415993
rect 442630 415919 442686 415928
rect 442078 343360 442134 343369
rect 442078 343295 442134 343304
rect 442184 341465 442212 415919
rect 442262 369200 442318 369209
rect 442262 369135 442264 369144
rect 442316 369135 442318 369144
rect 442264 369106 442316 369112
rect 442262 367024 442318 367033
rect 442262 366959 442318 366968
rect 442170 341456 442226 341465
rect 442170 341391 442226 341400
rect 441988 318844 442040 318850
rect 441988 318786 442040 318792
rect 441896 309120 441948 309126
rect 441896 309062 441948 309068
rect 441896 298104 441948 298110
rect 441896 298046 441948 298052
rect 441908 296070 441936 298046
rect 441896 296064 441948 296070
rect 441896 296006 441948 296012
rect 442000 286521 442028 318786
rect 442276 296886 442304 366959
rect 442446 365936 442502 365945
rect 442446 365871 442502 365880
rect 442460 298110 442488 365871
rect 443012 349897 443040 433327
rect 443104 431118 443132 431149
rect 443092 431112 443144 431118
rect 443090 431080 443092 431089
rect 443144 431080 443146 431089
rect 443090 431015 443146 431024
rect 442998 349888 443054 349897
rect 442998 349823 443054 349832
rect 443104 348809 443132 431015
rect 443288 418305 443316 486367
rect 443366 484800 443422 484809
rect 443366 484735 443422 484744
rect 443274 418296 443330 418305
rect 443274 418231 443330 418240
rect 443380 414905 443408 484735
rect 443472 447166 443500 488951
rect 443564 455462 443592 491302
rect 443552 455456 443604 455462
rect 443552 455398 443604 455404
rect 443460 447160 443512 447166
rect 443460 447102 443512 447108
rect 443656 437510 443684 495343
rect 443840 439113 443868 496431
rect 443920 491224 443972 491230
rect 443920 491166 443972 491172
rect 443932 490113 443960 491166
rect 443918 490104 443974 490113
rect 443918 490039 443974 490048
rect 443826 439104 443882 439113
rect 443826 439039 443882 439048
rect 443644 437504 443696 437510
rect 443644 437446 443696 437452
rect 443932 425241 443960 490039
rect 444392 460934 444420 512615
rect 444576 512145 444604 512722
rect 444562 512136 444618 512145
rect 444562 512071 444618 512080
rect 444392 460906 444512 460934
rect 444484 440366 444512 460906
rect 444472 440360 444524 440366
rect 444472 440302 444524 440308
rect 444194 439104 444250 439113
rect 444194 439039 444196 439048
rect 444248 439039 444250 439048
rect 444196 439010 444248 439016
rect 444380 437504 444432 437510
rect 444380 437446 444432 437452
rect 444392 436801 444420 437446
rect 444378 436792 444434 436801
rect 444378 436727 444380 436736
rect 444432 436727 444434 436736
rect 444380 436698 444432 436704
rect 444484 436642 444512 440302
rect 444392 436614 444512 436642
rect 443550 425232 443606 425241
rect 443550 425167 443606 425176
rect 443918 425232 443974 425241
rect 443918 425167 443974 425176
rect 443458 418296 443514 418305
rect 443458 418231 443514 418240
rect 443366 414896 443422 414905
rect 443366 414831 443422 414840
rect 443366 350568 443422 350577
rect 443366 350503 443422 350512
rect 443090 348800 443146 348809
rect 443090 348735 443146 348744
rect 443104 345014 443132 348735
rect 443276 347744 443328 347750
rect 443276 347686 443328 347692
rect 443104 344986 443224 345014
rect 442998 342816 443054 342825
rect 442998 342751 443054 342760
rect 442448 298104 442500 298110
rect 442448 298046 442500 298052
rect 442460 297634 442488 298046
rect 442448 297628 442500 297634
rect 442448 297570 442500 297576
rect 442264 296880 442316 296886
rect 442264 296822 442316 296828
rect 442276 296714 442304 296822
rect 442092 296686 442304 296714
rect 442092 296002 442120 296686
rect 442080 295996 442132 296002
rect 442080 295938 442132 295944
rect 441986 286512 442042 286521
rect 441986 286447 442042 286456
rect 441802 275768 441858 275777
rect 441802 275703 441858 275712
rect 443012 274417 443040 342751
rect 443090 341456 443146 341465
rect 443090 341391 443146 341400
rect 442998 274408 443054 274417
rect 442998 274343 443054 274352
rect 443104 272105 443132 341391
rect 443196 287201 443224 344986
rect 443288 318850 443316 347686
rect 443276 318844 443328 318850
rect 443276 318786 443328 318792
rect 443276 297492 443328 297498
rect 443276 297434 443328 297440
rect 443288 296546 443316 297434
rect 443276 296540 443328 296546
rect 443276 296482 443328 296488
rect 443380 291825 443408 350503
rect 443472 342825 443500 418231
rect 443564 346089 443592 425167
rect 443826 421832 443882 421841
rect 443826 421767 443882 421776
rect 443840 420918 443868 421767
rect 443828 420912 443880 420918
rect 443828 420854 443880 420860
rect 443840 412634 443868 420854
rect 444194 414896 444250 414905
rect 444194 414831 444196 414840
rect 444248 414831 444250 414840
rect 444196 414802 444248 414808
rect 443656 412606 443868 412634
rect 443550 346080 443606 346089
rect 443550 346015 443606 346024
rect 443656 344457 443684 412606
rect 444392 368665 444420 436614
rect 444470 434480 444526 434489
rect 444470 434415 444472 434424
rect 444524 434415 444526 434424
rect 444472 434386 444524 434392
rect 444472 432948 444524 432954
rect 444472 432890 444524 432896
rect 444484 432177 444512 432890
rect 444470 432168 444526 432177
rect 444470 432103 444526 432112
rect 444470 419520 444526 419529
rect 444470 419455 444472 419464
rect 444524 419455 444526 419464
rect 444472 419426 444524 419432
rect 444472 369912 444524 369918
rect 444472 369854 444524 369860
rect 444378 368656 444434 368665
rect 444378 368591 444434 368600
rect 444288 367056 444340 367062
rect 444288 366998 444340 367004
rect 444300 366489 444328 366998
rect 444286 366480 444342 366489
rect 444286 366415 444342 366424
rect 444194 365392 444250 365401
rect 444194 365327 444250 365336
rect 444208 364410 444236 365327
rect 444196 364404 444248 364410
rect 444196 364346 444248 364352
rect 443828 350532 443880 350538
rect 443828 350474 443880 350480
rect 443734 349888 443790 349897
rect 443734 349823 443790 349832
rect 443642 344448 443698 344457
rect 443642 344383 443698 344392
rect 443458 342816 443514 342825
rect 443458 342751 443514 342760
rect 443656 342310 443684 344383
rect 443644 342304 443696 342310
rect 443644 342246 443696 342252
rect 443644 326324 443696 326330
rect 443644 326266 443696 326272
rect 443656 296138 443684 326266
rect 443644 296132 443696 296138
rect 443644 296074 443696 296080
rect 443748 293026 443776 349823
rect 443564 292998 443776 293026
rect 443366 291816 443422 291825
rect 443366 291751 443422 291760
rect 443564 289513 443592 292998
rect 443642 292904 443698 292913
rect 443840 292890 443868 350474
rect 444208 326330 444236 364346
rect 444196 326324 444248 326330
rect 444196 326266 444248 326272
rect 444300 297498 444328 366415
rect 444484 362681 444512 369854
rect 444576 367878 444604 512071
rect 444746 510504 444802 510513
rect 444746 510439 444802 510448
rect 444656 499520 444708 499526
rect 444656 499462 444708 499468
rect 444668 498681 444696 499462
rect 444654 498672 444710 498681
rect 444654 498607 444710 498616
rect 444656 493332 444708 493338
rect 444656 493274 444708 493280
rect 444668 492833 444696 493274
rect 444654 492824 444710 492833
rect 444654 492759 444710 492768
rect 444654 487928 444710 487937
rect 444654 487863 444656 487872
rect 444708 487863 444710 487872
rect 444656 487834 444708 487840
rect 444654 484256 444710 484265
rect 444654 484191 444656 484200
rect 444708 484191 444710 484200
rect 444656 484162 444708 484168
rect 444654 438016 444710 438025
rect 444654 437951 444656 437960
rect 444708 437951 444710 437960
rect 444656 437922 444708 437928
rect 444654 417208 444710 417217
rect 444654 417143 444656 417152
rect 444708 417143 444710 417152
rect 444656 417114 444708 417120
rect 444564 367872 444616 367878
rect 444564 367814 444616 367820
rect 444760 367062 444788 510439
rect 444852 369209 444880 513159
rect 444944 369753 444972 513742
rect 445392 512644 445444 512650
rect 445392 512586 445444 512592
rect 445404 511057 445432 512586
rect 445668 511964 445720 511970
rect 445668 511906 445720 511912
rect 445680 511601 445708 511906
rect 445666 511592 445722 511601
rect 445666 511527 445722 511536
rect 445390 511048 445446 511057
rect 445390 510983 445446 510992
rect 445298 504112 445354 504121
rect 445298 504047 445354 504056
rect 445312 503742 445340 504047
rect 445300 503736 445352 503742
rect 445300 503678 445352 503684
rect 445114 503568 445170 503577
rect 445114 503503 445170 503512
rect 445022 503024 445078 503033
rect 445022 502959 445078 502968
rect 445036 460222 445064 502959
rect 445128 499574 445156 503503
rect 445206 502480 445262 502489
rect 445206 502415 445262 502424
rect 445220 502314 445248 502415
rect 445208 502308 445260 502314
rect 445208 502250 445260 502256
rect 445220 500834 445248 502250
rect 445298 501392 445354 501401
rect 445298 501327 445354 501336
rect 445312 501022 445340 501327
rect 445300 501016 445352 501022
rect 445300 500958 445352 500964
rect 445220 500806 445340 500834
rect 445128 499546 445248 499574
rect 445116 485784 445168 485790
rect 445114 485752 445116 485761
rect 445168 485752 445170 485761
rect 445114 485687 445170 485696
rect 445024 460216 445076 460222
rect 445024 460158 445076 460164
rect 444930 369744 444986 369753
rect 444930 369679 444986 369688
rect 444838 369200 444894 369209
rect 444838 369135 444894 369144
rect 444748 367056 444800 367062
rect 444748 366998 444800 367004
rect 444654 365936 444710 365945
rect 444654 365871 444710 365880
rect 444668 365770 444696 365871
rect 444656 365764 444708 365770
rect 444656 365706 444708 365712
rect 444932 365696 444984 365702
rect 444932 365638 444984 365644
rect 444944 364857 444972 365638
rect 444930 364848 444986 364857
rect 444930 364783 444986 364792
rect 444470 362672 444526 362681
rect 444470 362607 444526 362616
rect 445036 359009 445064 460158
rect 445220 441726 445248 499546
rect 445312 494766 445340 500806
rect 445300 494760 445352 494766
rect 445300 494702 445352 494708
rect 445300 494624 445352 494630
rect 445300 494566 445352 494572
rect 445312 494329 445340 494566
rect 445298 494320 445354 494329
rect 445298 494255 445354 494264
rect 445300 493400 445352 493406
rect 445298 493368 445300 493377
rect 445352 493368 445354 493377
rect 445298 493303 445354 493312
rect 445298 491192 445354 491201
rect 445298 491127 445354 491136
rect 445312 491094 445340 491127
rect 445300 491088 445352 491094
rect 445300 491030 445352 491036
rect 445298 487384 445354 487393
rect 445298 487319 445300 487328
rect 445352 487319 445354 487328
rect 445300 487290 445352 487296
rect 445300 442944 445352 442950
rect 445300 442886 445352 442892
rect 445312 441794 445340 442886
rect 445300 441788 445352 441794
rect 445300 441730 445352 441736
rect 445208 441720 445260 441726
rect 445208 441662 445260 441668
rect 445114 441416 445170 441425
rect 445114 441351 445116 441360
rect 445168 441351 445170 441360
rect 445116 441322 445168 441328
rect 445116 436824 445168 436830
rect 445116 436766 445168 436772
rect 445128 364018 445156 436766
rect 445220 364334 445248 441662
rect 445312 436830 445340 441730
rect 445300 436824 445352 436830
rect 445300 436766 445352 436772
rect 445404 367033 445432 510983
rect 445668 509992 445720 509998
rect 445666 509960 445668 509969
rect 445720 509960 445722 509969
rect 445576 509924 445628 509930
rect 445666 509895 445722 509904
rect 445576 509866 445628 509872
rect 445588 509425 445616 509866
rect 445574 509416 445630 509425
rect 445574 509351 445630 509360
rect 445574 508872 445630 508881
rect 445574 508807 445630 508816
rect 445588 507890 445616 508807
rect 445668 508564 445720 508570
rect 445668 508506 445720 508512
rect 445680 508337 445708 508506
rect 445666 508328 445722 508337
rect 445666 508263 445722 508272
rect 445576 507884 445628 507890
rect 445576 507826 445628 507832
rect 445574 507240 445630 507249
rect 445574 507175 445576 507184
rect 445628 507175 445630 507184
rect 445576 507146 445628 507152
rect 445668 507136 445720 507142
rect 445668 507078 445720 507084
rect 445680 506705 445708 507078
rect 445666 506696 445722 506705
rect 445666 506631 445722 506640
rect 445666 506152 445722 506161
rect 445666 506087 445722 506096
rect 445576 505912 445628 505918
rect 445576 505854 445628 505860
rect 445588 505617 445616 505854
rect 445574 505608 445630 505617
rect 445574 505543 445630 505552
rect 445680 505170 445708 506087
rect 445668 505164 445720 505170
rect 445668 505106 445720 505112
rect 445666 504520 445722 504529
rect 445666 504455 445722 504464
rect 445680 504422 445708 504455
rect 445668 504416 445720 504422
rect 445668 504358 445720 504364
rect 445482 501936 445538 501945
rect 445482 501871 445538 501880
rect 445496 500954 445524 501871
rect 445484 500948 445536 500954
rect 445484 500890 445536 500896
rect 445496 499574 445524 500890
rect 445576 500880 445628 500886
rect 445576 500822 445628 500828
rect 445588 500313 445616 500822
rect 445668 500812 445720 500818
rect 445668 500754 445720 500760
rect 445574 500304 445630 500313
rect 445574 500239 445630 500248
rect 445680 499769 445708 500754
rect 445666 499760 445722 499769
rect 445666 499695 445722 499704
rect 445496 499546 445708 499574
rect 445574 499216 445630 499225
rect 445574 499151 445630 499160
rect 445588 498234 445616 499151
rect 445576 498228 445628 498234
rect 445576 498170 445628 498176
rect 445482 498128 445538 498137
rect 445482 498063 445538 498072
rect 445496 497826 445524 498063
rect 445484 497820 445536 497826
rect 445484 497762 445536 497768
rect 445574 497040 445630 497049
rect 445574 496975 445576 496984
rect 445628 496975 445630 496984
rect 445576 496946 445628 496952
rect 445576 494760 445628 494766
rect 445576 494702 445628 494708
rect 445482 488472 445538 488481
rect 445482 488407 445538 488416
rect 445496 487218 445524 488407
rect 445484 487212 445536 487218
rect 445484 487154 445536 487160
rect 445482 486296 445538 486305
rect 445482 486231 445538 486240
rect 445496 485858 445524 486231
rect 445484 485852 445536 485858
rect 445484 485794 445536 485800
rect 445482 484664 445538 484673
rect 445482 484599 445484 484608
rect 445536 484599 445538 484608
rect 445484 484570 445536 484576
rect 445588 442950 445616 494702
rect 445576 442944 445628 442950
rect 445576 442886 445628 442892
rect 445574 440328 445630 440337
rect 445574 440263 445576 440272
rect 445628 440263 445630 440272
rect 445576 440234 445628 440240
rect 445576 426896 445628 426902
rect 445576 426838 445628 426844
rect 445588 426465 445616 426838
rect 445574 426456 445630 426465
rect 445574 426391 445630 426400
rect 445576 420640 445628 420646
rect 445574 420608 445576 420617
rect 445628 420608 445630 420617
rect 445574 420543 445630 420552
rect 445484 413704 445536 413710
rect 445482 413672 445484 413681
rect 445536 413672 445538 413681
rect 445482 413607 445538 413616
rect 445484 412616 445536 412622
rect 445482 412584 445484 412593
rect 445536 412584 445538 412593
rect 445482 412519 445538 412528
rect 445390 367024 445446 367033
rect 445390 366959 445446 366968
rect 445576 364336 445628 364342
rect 445220 364306 445340 364334
rect 445128 363990 445248 364018
rect 445116 363860 445168 363866
rect 445116 363802 445168 363808
rect 445128 363225 445156 363802
rect 445114 363216 445170 363225
rect 445114 363151 445170 363160
rect 445116 362908 445168 362914
rect 445116 362850 445168 362856
rect 445128 362137 445156 362850
rect 445114 362128 445170 362137
rect 445114 362063 445170 362072
rect 445114 361584 445170 361593
rect 445114 361519 445116 361528
rect 445168 361519 445170 361528
rect 445116 361490 445168 361496
rect 445114 360496 445170 360505
rect 445114 360431 445170 360440
rect 445128 360194 445156 360431
rect 445116 360188 445168 360194
rect 445116 360130 445168 360136
rect 445114 359544 445170 359553
rect 445114 359479 445170 359488
rect 445022 359000 445078 359009
rect 444944 358958 445022 358986
rect 444746 358456 444802 358465
rect 444746 358391 444802 358400
rect 444654 354648 444710 354657
rect 444654 354583 444710 354592
rect 444668 353326 444696 354583
rect 444656 353320 444708 353326
rect 444656 353262 444708 353268
rect 444380 351416 444432 351422
rect 444378 351384 444380 351393
rect 444432 351384 444434 351393
rect 444378 351319 444434 351328
rect 444392 350538 444420 351319
rect 444380 350532 444432 350538
rect 444380 350474 444432 350480
rect 444378 347712 444434 347721
rect 444378 347647 444434 347656
rect 444392 346730 444420 347647
rect 444380 346724 444432 346730
rect 444380 346666 444432 346672
rect 444470 344992 444526 345001
rect 444470 344927 444526 344936
rect 444380 343936 444432 343942
rect 444378 343904 444380 343913
rect 444432 343904 444434 343913
rect 444378 343839 444434 343848
rect 444380 297560 444432 297566
rect 444378 297528 444380 297537
rect 444432 297528 444434 297537
rect 444288 297492 444340 297498
rect 444378 297463 444434 297472
rect 444288 297434 444340 297440
rect 444300 296954 444328 297434
rect 444288 296948 444340 296954
rect 444288 296890 444340 296896
rect 444380 296540 444432 296546
rect 444380 296482 444432 296488
rect 444392 296449 444420 296482
rect 444378 296440 444434 296449
rect 444378 296375 444434 296384
rect 443698 292862 443868 292890
rect 443642 292839 443698 292848
rect 443550 289504 443606 289513
rect 443550 289439 443606 289448
rect 443182 287192 443238 287201
rect 443182 287127 443184 287136
rect 443236 287127 443238 287136
rect 443184 287098 443236 287104
rect 443196 287067 443224 287098
rect 443090 272096 443146 272105
rect 443090 272031 443146 272040
rect 441618 271552 441674 271561
rect 441618 271487 441674 271496
rect 441632 270094 441660 271487
rect 441620 270088 441672 270094
rect 441620 270030 441672 270036
rect 440956 268668 441108 268682
rect 440942 268654 441108 268668
rect 440942 268546 440970 268654
rect 432524 268532 432952 268546
rect 440620 268532 440970 268546
rect 432524 268518 432966 268532
rect 432938 267866 432966 268518
rect 440620 268518 440956 268532
rect 434884 268110 434944 268138
rect 436908 268110 436968 268138
rect 432892 267838 432966 267866
rect 431868 266280 431920 266286
rect 431868 266222 431920 266228
rect 432892 265742 432920 267838
rect 434916 266354 434944 268110
rect 434904 266348 434956 266354
rect 434904 266290 434956 266296
rect 431960 265736 432012 265742
rect 431960 265678 432012 265684
rect 432880 265736 432932 265742
rect 432880 265678 432932 265684
rect 431972 209774 432000 265678
rect 434916 265033 434944 266290
rect 436940 266286 436968 268110
rect 438918 268002 438946 268124
rect 438872 267974 438946 268002
rect 436928 266280 436980 266286
rect 436928 266222 436980 266228
rect 436940 265577 436968 266222
rect 438872 266218 438900 267974
rect 438860 266212 438912 266218
rect 438860 266154 438912 266160
rect 440620 265674 440648 268518
rect 440608 265668 440660 265674
rect 440608 265610 440660 265616
rect 441068 265668 441120 265674
rect 441068 265610 441120 265616
rect 436926 265568 436982 265577
rect 436926 265503 436982 265512
rect 434902 265024 434958 265033
rect 434902 264959 434958 264968
rect 431972 209746 432552 209774
rect 432524 196058 432552 209746
rect 435178 196072 435234 196081
rect 432524 196030 432952 196058
rect 434732 196030 435178 196058
rect 432524 180794 432552 196030
rect 431972 180766 432552 180794
rect 431868 153876 431920 153882
rect 431868 153818 431920 153824
rect 431316 153332 431368 153338
rect 431316 153274 431368 153280
rect 431328 142118 431356 153274
rect 431408 151972 431460 151978
rect 431408 151914 431460 151920
rect 431420 143546 431448 151914
rect 431408 143540 431460 143546
rect 431408 143482 431460 143488
rect 431316 142112 431368 142118
rect 431316 142054 431368 142060
rect 431316 138780 431368 138786
rect 431316 138722 431368 138728
rect 431328 124166 431356 138722
rect 431316 124160 431368 124166
rect 431316 124102 431368 124108
rect 431880 122806 431908 153818
rect 431972 132494 432000 180766
rect 434732 153882 434760 196030
rect 435178 196007 435234 196016
rect 436742 196072 436798 196081
rect 441080 196058 441108 265610
rect 442080 258732 442132 258738
rect 442080 258674 442132 258680
rect 441712 255332 441764 255338
rect 441712 255274 441764 255280
rect 441620 226296 441672 226302
rect 441618 226264 441620 226273
rect 441672 226264 441674 226273
rect 441618 226199 441674 226208
rect 441620 226160 441672 226166
rect 441620 226102 441672 226108
rect 441632 225593 441660 226102
rect 441618 225584 441674 225593
rect 441618 225519 441674 225528
rect 441724 225026 441752 255274
rect 441804 251252 441856 251258
rect 441804 251194 441856 251200
rect 441816 228342 441844 251194
rect 441896 249076 441948 249082
rect 441896 249018 441948 249024
rect 441804 228336 441856 228342
rect 441804 228278 441856 228284
rect 441908 225146 441936 249018
rect 441988 246356 442040 246362
rect 441988 246298 442040 246304
rect 442000 225214 442028 246298
rect 441988 225208 442040 225214
rect 441988 225150 442040 225156
rect 441896 225140 441948 225146
rect 441896 225082 441948 225088
rect 441724 224998 442028 225026
rect 441712 224936 441764 224942
rect 441618 224904 441674 224913
rect 441712 224878 441764 224884
rect 441618 224839 441620 224848
rect 441672 224839 441674 224848
rect 441620 224810 441672 224816
rect 441724 224505 441752 224878
rect 441710 224496 441766 224505
rect 441710 224431 441766 224440
rect 441804 223916 441856 223922
rect 441804 223858 441856 223864
rect 441816 220697 441844 223858
rect 442000 223417 442028 224998
rect 442092 223553 442120 258674
rect 443104 258074 443132 272031
rect 443012 258046 443132 258074
rect 442356 228336 442408 228342
rect 442356 228278 442408 228284
rect 442264 225208 442316 225214
rect 442264 225150 442316 225156
rect 442172 225140 442224 225146
rect 442172 225082 442224 225088
rect 442078 223544 442134 223553
rect 442078 223479 442134 223488
rect 441986 223408 442042 223417
rect 441986 223343 442042 223352
rect 442184 221921 442212 225082
rect 442170 221912 442226 221921
rect 442170 221847 442226 221856
rect 442276 221377 442304 225150
rect 442368 222465 442396 228278
rect 442354 222456 442410 222465
rect 442354 222391 442410 222400
rect 442262 221368 442318 221377
rect 442262 221303 442318 221312
rect 441802 220688 441858 220697
rect 441802 220623 441858 220632
rect 442724 212424 442776 212430
rect 442724 212366 442776 212372
rect 442736 211721 442764 212366
rect 442262 211712 442318 211721
rect 442262 211647 442318 211656
rect 442722 211712 442778 211721
rect 442722 211647 442778 211656
rect 442172 211064 442224 211070
rect 442172 211006 442224 211012
rect 442184 210633 442212 211006
rect 442170 210624 442226 210633
rect 442170 210559 442226 210568
rect 442078 205864 442134 205873
rect 442078 205799 442134 205808
rect 441618 205048 441674 205057
rect 441618 204983 441674 204992
rect 436798 196030 437336 196058
rect 438932 196030 438992 196058
rect 440956 196030 441108 196058
rect 436742 196007 436798 196016
rect 437308 190454 437336 196030
rect 438964 193866 438992 196030
rect 438952 193860 439004 193866
rect 438952 193802 439004 193808
rect 437308 190426 437428 190454
rect 437400 154222 437428 190426
rect 437388 154216 437440 154222
rect 437388 154158 437440 154164
rect 434720 153876 434772 153882
rect 434720 153818 434772 153824
rect 431972 132466 432552 132494
rect 432524 124794 432552 132466
rect 441080 124794 441108 196030
rect 441632 155378 441660 204983
rect 441802 204640 441858 204649
rect 441802 204575 441858 204584
rect 441710 201920 441766 201929
rect 441710 201855 441766 201864
rect 441724 166994 441752 201855
rect 441816 168366 441844 204575
rect 441986 203552 442042 203561
rect 441986 203487 442042 203496
rect 442000 176662 442028 203487
rect 442092 180794 442120 205799
rect 442184 184210 442212 210559
rect 442276 191146 442304 211647
rect 442908 205352 442960 205358
rect 442906 205320 442908 205329
rect 442960 205320 442962 205329
rect 442906 205255 442962 205264
rect 442724 203992 442776 203998
rect 442724 203934 442776 203940
rect 442736 203697 442764 203934
rect 442722 203688 442778 203697
rect 442722 203623 442778 203632
rect 442356 203380 442408 203386
rect 442356 203322 442408 203328
rect 442368 203153 442396 203322
rect 442354 203144 442410 203153
rect 442354 203079 442410 203088
rect 442368 200114 442396 203079
rect 442908 202768 442960 202774
rect 442908 202710 442960 202716
rect 442920 202065 442948 202710
rect 442906 202056 442962 202065
rect 442906 201991 442962 202000
rect 442368 200086 442488 200114
rect 442264 191140 442316 191146
rect 442264 191082 442316 191088
rect 442172 184204 442224 184210
rect 442172 184146 442224 184152
rect 442092 180766 442304 180794
rect 442276 178702 442304 180766
rect 442264 178696 442316 178702
rect 442264 178638 442316 178644
rect 441988 176656 442040 176662
rect 441988 176598 442040 176604
rect 442000 175302 442028 176598
rect 441988 175296 442040 175302
rect 441988 175238 442040 175244
rect 441804 168360 441856 168366
rect 441804 168302 441856 168308
rect 441724 166966 441936 166994
rect 441908 165578 441936 166966
rect 441896 165572 441948 165578
rect 441896 165514 441948 165520
rect 441620 155372 441672 155378
rect 441620 155314 441672 155320
rect 441632 154358 441660 155314
rect 441804 154556 441856 154562
rect 441804 154498 441856 154504
rect 441620 154352 441672 154358
rect 441620 154294 441672 154300
rect 441712 154216 441764 154222
rect 441712 154158 441764 154164
rect 441618 135960 441674 135969
rect 441618 135895 441620 135904
rect 441672 135895 441674 135904
rect 441620 135866 441672 135872
rect 441632 125322 441660 135866
rect 441620 125316 441672 125322
rect 441620 125258 441672 125264
rect 441618 124944 441674 124953
rect 441618 124879 441620 124888
rect 441672 124879 441674 124888
rect 441620 124850 441672 124856
rect 432524 124766 433012 124794
rect 440956 124766 441292 124794
rect 432984 124522 433012 124766
rect 432984 124494 433196 124522
rect 431868 122800 431920 122806
rect 431868 122742 431920 122748
rect 433168 122738 433196 124494
rect 434732 124086 434884 124114
rect 436908 124086 437244 124114
rect 434732 122806 434760 124086
rect 434720 122800 434772 122806
rect 434720 122742 434772 122748
rect 433156 122732 433208 122738
rect 433156 122674 433208 122680
rect 437216 122670 437244 124086
rect 438918 123842 438946 124100
rect 438872 123814 438946 123842
rect 437204 122664 437256 122670
rect 437204 122606 437256 122612
rect 438872 122602 438900 123814
rect 441264 122806 441292 124766
rect 441252 122800 441304 122806
rect 441252 122742 441304 122748
rect 441724 122670 441752 154158
rect 441816 154057 441844 154498
rect 441802 154048 441858 154057
rect 441802 153983 441858 153992
rect 442276 153542 442304 178638
rect 442356 175296 442408 175302
rect 442356 175238 442408 175244
rect 442368 154426 442396 175238
rect 442460 171834 442488 200086
rect 443012 197713 443040 258046
rect 443552 242956 443604 242962
rect 443552 242898 443604 242904
rect 443184 236700 443236 236706
rect 443184 236642 443236 236648
rect 443196 229094 443224 236642
rect 443276 233912 443328 233918
rect 443276 233854 443328 233860
rect 443104 229066 443224 229094
rect 443104 219745 443132 229066
rect 443184 224256 443236 224262
rect 443184 224198 443236 224204
rect 443090 219736 443146 219745
rect 443090 219671 443146 219680
rect 443196 219434 443224 224198
rect 443288 219570 443316 233854
rect 443368 231124 443420 231130
rect 443368 231066 443420 231072
rect 443276 219564 443328 219570
rect 443276 219506 443328 219512
rect 443196 219406 443316 219434
rect 443288 217569 443316 219406
rect 443380 218657 443408 231066
rect 443460 226364 443512 226370
rect 443460 226306 443512 226312
rect 443366 218648 443422 218657
rect 443366 218583 443422 218592
rect 443380 218074 443408 218583
rect 443472 218113 443500 226306
rect 443564 220833 443592 242898
rect 443656 238406 443684 292839
rect 444288 289876 444340 289882
rect 444288 289818 444340 289824
rect 444300 289513 444328 289818
rect 444286 289504 444342 289513
rect 444286 289439 444342 289448
rect 444380 282872 444432 282878
rect 444380 282814 444432 282820
rect 444392 282577 444420 282814
rect 444378 282568 444434 282577
rect 444378 282503 444434 282512
rect 444484 280129 444512 344927
rect 444656 342304 444708 342310
rect 444656 342246 444708 342252
rect 444562 340232 444618 340241
rect 444562 340167 444618 340176
rect 444576 339522 444604 340167
rect 444564 339516 444616 339522
rect 444564 339458 444616 339464
rect 444564 309120 444616 309126
rect 444564 309062 444616 309068
rect 444470 280120 444526 280129
rect 444470 280055 444526 280064
rect 444576 276729 444604 309062
rect 444668 277953 444696 342246
rect 444760 297090 444788 358391
rect 444944 297158 444972 358958
rect 445022 358935 445078 358944
rect 445022 355736 445078 355745
rect 445022 355671 445078 355680
rect 445036 355366 445064 355671
rect 445024 355360 445076 355366
rect 445024 355302 445076 355308
rect 444932 297152 444984 297158
rect 444932 297094 444984 297100
rect 444748 297084 444800 297090
rect 444748 297026 444800 297032
rect 444760 296714 444788 297026
rect 444760 296686 444880 296714
rect 444746 284880 444802 284889
rect 444746 284815 444748 284824
rect 444800 284815 444802 284824
rect 444748 284786 444800 284792
rect 444746 281344 444802 281353
rect 444746 281279 444748 281288
rect 444800 281279 444802 281288
rect 444748 281250 444800 281256
rect 444654 277944 444710 277953
rect 444654 277879 444710 277888
rect 444562 276720 444618 276729
rect 444562 276655 444618 276664
rect 444562 273320 444618 273329
rect 444562 273255 444618 273264
rect 444576 273222 444604 273255
rect 444564 273216 444616 273222
rect 444564 273158 444616 273164
rect 444576 268394 444604 273158
rect 444564 268388 444616 268394
rect 444564 268330 444616 268336
rect 444380 247920 444432 247926
rect 444380 247862 444432 247868
rect 444392 247722 444420 247862
rect 444380 247716 444432 247722
rect 444380 247658 444432 247664
rect 443644 238400 443696 238406
rect 443644 238342 443696 238348
rect 444288 238400 444340 238406
rect 444288 238342 444340 238348
rect 444300 238066 444328 238342
rect 444288 238060 444340 238066
rect 444288 238002 444340 238008
rect 443550 220824 443606 220833
rect 443550 220759 443606 220768
rect 443644 219428 443696 219434
rect 443644 219370 443696 219376
rect 443656 219201 443684 219370
rect 443642 219192 443698 219201
rect 443642 219127 443698 219136
rect 443656 218142 443684 219127
rect 443644 218136 443696 218142
rect 443458 218104 443514 218113
rect 443368 218068 443420 218074
rect 443644 218078 443696 218084
rect 443458 218039 443514 218048
rect 443368 218010 443420 218016
rect 443274 217560 443330 217569
rect 443274 217495 443330 217504
rect 443288 216714 443316 217495
rect 443276 216708 443328 216714
rect 443276 216650 443328 216656
rect 443366 212800 443422 212809
rect 443366 212735 443422 212744
rect 443274 212256 443330 212265
rect 443274 212191 443330 212200
rect 443184 211132 443236 211138
rect 443184 211074 443236 211080
rect 443196 210089 443224 211074
rect 443182 210080 443238 210089
rect 443182 210015 443238 210024
rect 443196 200114 443224 210015
rect 443104 200086 443224 200114
rect 442998 197704 443054 197713
rect 442998 197639 443054 197648
rect 443104 181490 443132 200086
rect 443288 194478 443316 212191
rect 443380 197266 443408 212735
rect 443458 211168 443514 211177
rect 443458 211103 443514 211112
rect 443368 197260 443420 197266
rect 443368 197202 443420 197208
rect 443276 194472 443328 194478
rect 443276 194414 443328 194420
rect 443472 187678 443500 211103
rect 444300 207369 444328 238002
rect 444392 215529 444420 247658
rect 444472 242888 444524 242894
rect 444472 242830 444524 242836
rect 444484 224618 444512 242830
rect 444564 241460 444616 241466
rect 444564 241402 444616 241408
rect 444576 240174 444604 241402
rect 444564 240168 444616 240174
rect 444564 240110 444616 240116
rect 444576 229094 444604 240110
rect 444668 240106 444696 277879
rect 444746 274408 444802 274417
rect 444746 274343 444802 274352
rect 444656 240100 444708 240106
rect 444656 240042 444708 240048
rect 444760 238754 444788 274343
rect 444852 241466 444880 296686
rect 444944 242894 444972 297094
rect 444932 242888 444984 242894
rect 444932 242830 444984 242836
rect 444840 241460 444892 241466
rect 444840 241402 444892 241408
rect 444760 238726 444972 238754
rect 444944 231130 444972 238726
rect 444932 231124 444984 231130
rect 444932 231066 444984 231072
rect 444840 230444 444892 230450
rect 444840 230386 444892 230392
rect 444852 229770 444880 230386
rect 444840 229764 444892 229770
rect 444840 229706 444892 229712
rect 444576 229066 444696 229094
rect 444484 224590 444604 224618
rect 444472 224324 444524 224330
rect 444472 224266 444524 224272
rect 444484 216073 444512 224266
rect 444470 216064 444526 216073
rect 444470 215999 444526 216008
rect 444484 215898 444512 215999
rect 444472 215892 444524 215898
rect 444472 215834 444524 215840
rect 444378 215520 444434 215529
rect 444378 215455 444434 215464
rect 444576 214985 444604 224590
rect 444562 214976 444618 214985
rect 444562 214911 444618 214920
rect 444668 214441 444696 229066
rect 444746 223544 444802 223553
rect 444746 223479 444802 223488
rect 444760 222358 444788 223479
rect 444748 222352 444800 222358
rect 444748 222294 444800 222300
rect 444746 221912 444802 221921
rect 444746 221847 444802 221856
rect 444760 220930 444788 221847
rect 444748 220924 444800 220930
rect 444748 220866 444800 220872
rect 444746 220280 444802 220289
rect 444746 220215 444802 220224
rect 444760 219570 444788 220215
rect 444748 219564 444800 219570
rect 444748 219506 444800 219512
rect 444654 214432 444710 214441
rect 444654 214367 444710 214376
rect 444852 213897 444880 229706
rect 444838 213888 444894 213897
rect 444838 213823 444894 213832
rect 444748 212492 444800 212498
rect 444748 212434 444800 212440
rect 444760 212265 444788 212434
rect 444746 212256 444802 212265
rect 444746 212191 444802 212200
rect 444564 209092 444616 209098
rect 444564 209034 444616 209040
rect 444286 207360 444342 207369
rect 444286 207295 444342 207304
rect 444194 206272 444250 206281
rect 444194 206207 444250 206216
rect 444208 205630 444236 206207
rect 444300 205766 444328 207295
rect 444380 205896 444432 205902
rect 444378 205864 444380 205873
rect 444432 205864 444434 205873
rect 444378 205799 444434 205808
rect 444288 205760 444340 205766
rect 444288 205702 444340 205708
rect 443644 205624 443696 205630
rect 443644 205566 443696 205572
rect 444196 205624 444248 205630
rect 444196 205566 444248 205572
rect 443460 187672 443512 187678
rect 443460 187614 443512 187620
rect 443092 181484 443144 181490
rect 443092 181426 443144 181432
rect 442724 172576 442776 172582
rect 442724 172518 442776 172524
rect 442448 171828 442500 171834
rect 442448 171770 442500 171776
rect 442460 154494 442488 171770
rect 442632 171080 442684 171086
rect 442632 171022 442684 171028
rect 442644 170406 442672 171022
rect 442632 170400 442684 170406
rect 442632 170342 442684 170348
rect 442448 154488 442500 154494
rect 442448 154430 442500 154436
rect 442356 154420 442408 154426
rect 442356 154362 442408 154368
rect 442264 153536 442316 153542
rect 442264 153478 442316 153484
rect 441804 152040 441856 152046
rect 441802 152008 441804 152017
rect 441856 152008 441858 152017
rect 441802 151943 441858 151952
rect 442276 146033 442304 153478
rect 442644 151842 442672 170342
rect 442736 152114 442764 172518
rect 443000 165572 443052 165578
rect 443000 165514 443052 165520
rect 442908 162852 442960 162858
rect 442908 162794 442960 162800
rect 442920 161498 442948 162794
rect 442908 161492 442960 161498
rect 442908 161434 442960 161440
rect 442814 158808 442870 158817
rect 442814 158743 442870 158752
rect 442724 152108 442776 152114
rect 442724 152050 442776 152056
rect 442632 151836 442684 151842
rect 442632 151778 442684 151784
rect 442736 150385 442764 152050
rect 442722 150376 442778 150385
rect 442722 150311 442778 150320
rect 442262 146024 442318 146033
rect 442262 145959 442318 145968
rect 442828 132530 442856 158743
rect 442920 133958 442948 161434
rect 443012 137329 443040 165514
rect 443656 158030 443684 205566
rect 444380 204808 444432 204814
rect 444378 204776 444380 204785
rect 444432 204776 444434 204785
rect 444378 204711 444434 204720
rect 444470 198792 444526 198801
rect 444470 198727 444526 198736
rect 443092 158024 443144 158030
rect 443092 157966 443144 157972
rect 443644 158024 443696 158030
rect 443644 157966 443696 157972
rect 443104 153406 443132 157966
rect 443092 153400 443144 153406
rect 443092 153342 443144 153348
rect 443104 146577 443132 153342
rect 444196 151836 444248 151842
rect 444196 151778 444248 151784
rect 444208 151722 444236 151778
rect 444208 151706 444420 151722
rect 444208 151700 444432 151706
rect 444208 151694 444380 151700
rect 444380 151642 444432 151648
rect 444392 147801 444420 151642
rect 444378 147792 444434 147801
rect 444378 147727 444434 147736
rect 443090 146568 443146 146577
rect 443090 146503 443146 146512
rect 442998 137320 443054 137329
rect 442998 137255 443054 137264
rect 443090 135008 443146 135017
rect 443090 134943 443146 134952
rect 443104 134026 443132 134943
rect 443092 134020 443144 134026
rect 443092 133962 443144 133968
rect 442908 133952 442960 133958
rect 442908 133894 442960 133900
rect 442816 132524 442868 132530
rect 442816 132466 442868 132472
rect 442906 129840 442962 129849
rect 442906 129775 442962 129784
rect 442920 127702 442948 129775
rect 442908 127696 442960 127702
rect 442908 127638 442960 127644
rect 441894 127528 441950 127537
rect 441894 127463 441950 127472
rect 441802 126440 441858 126449
rect 441802 126375 441858 126384
rect 441816 125526 441844 126375
rect 441908 126070 441936 127463
rect 441896 126064 441948 126070
rect 441896 126006 441948 126012
rect 442920 126002 442948 127638
rect 442908 125996 442960 126002
rect 442908 125938 442960 125944
rect 442078 125760 442134 125769
rect 442078 125695 442134 125704
rect 441804 125520 441856 125526
rect 441804 125462 441856 125468
rect 442092 125390 442120 125695
rect 443104 125458 443132 133962
rect 444196 132524 444248 132530
rect 444196 132466 444248 132472
rect 444208 132161 444236 132466
rect 444194 132152 444250 132161
rect 444194 132087 444250 132096
rect 444484 129849 444512 198727
rect 444576 154562 444604 209034
rect 444746 207904 444802 207913
rect 444746 207839 444802 207848
rect 444656 205760 444708 205766
rect 444656 205702 444708 205708
rect 444668 163810 444696 205702
rect 444760 172582 444788 207839
rect 444838 201376 444894 201385
rect 444838 201311 444894 201320
rect 444852 200433 444880 201311
rect 444838 200424 444894 200433
rect 444838 200359 444894 200368
rect 444748 172576 444800 172582
rect 444748 172518 444800 172524
rect 444852 167686 444880 200359
rect 444944 198801 444972 231066
rect 445036 212430 445064 355302
rect 445128 354674 445156 359479
rect 445220 358465 445248 363990
rect 445312 359553 445340 364306
rect 445574 364304 445576 364313
rect 445628 364304 445630 364313
rect 445574 364239 445630 364248
rect 445390 360088 445446 360097
rect 445390 360023 445446 360032
rect 445298 359544 445354 359553
rect 445298 359479 445354 359488
rect 445206 358456 445262 358465
rect 445206 358391 445262 358400
rect 445298 357368 445354 357377
rect 445298 357303 445354 357312
rect 445128 354646 445248 354674
rect 445116 353864 445168 353870
rect 445116 353806 445168 353812
rect 445128 353569 445156 353806
rect 445114 353560 445170 353569
rect 445114 353495 445170 353504
rect 445116 346656 445168 346662
rect 445114 346624 445116 346633
rect 445168 346624 445170 346633
rect 445114 346559 445170 346568
rect 445116 342304 445168 342310
rect 445114 342272 445116 342281
rect 445168 342272 445170 342281
rect 445114 342207 445170 342216
rect 445116 298036 445168 298042
rect 445116 297978 445168 297984
rect 445128 297226 445156 297978
rect 445116 297220 445168 297226
rect 445116 297162 445168 297168
rect 445128 230450 445156 297162
rect 445220 296002 445248 354646
rect 445312 298110 445340 357303
rect 445300 298104 445352 298110
rect 445300 298046 445352 298052
rect 445404 297294 445432 360023
rect 445680 358766 445708 499546
rect 445772 497593 445800 585398
rect 446404 585336 446456 585342
rect 446404 585278 446456 585284
rect 445850 582040 445906 582049
rect 445850 581975 445906 581984
rect 445758 497584 445814 497593
rect 445758 497519 445814 497528
rect 445772 496874 445800 497519
rect 445760 496868 445812 496874
rect 445760 496810 445812 496816
rect 445864 495961 445892 581975
rect 445942 572792 445998 572801
rect 445942 572727 445998 572736
rect 445850 495952 445906 495961
rect 445850 495887 445906 495896
rect 445864 491178 445892 495887
rect 445956 491298 445984 572727
rect 446416 513806 446444 585278
rect 447784 583908 447836 583914
rect 447784 583850 447836 583856
rect 446496 564596 446548 564602
rect 446496 564538 446548 564544
rect 446508 523734 446536 564538
rect 446588 561196 446640 561202
rect 446588 561138 446640 561144
rect 446496 523728 446548 523734
rect 446496 523670 446548 523676
rect 446404 513800 446456 513806
rect 446404 513742 446456 513748
rect 446404 503668 446456 503674
rect 446404 503610 446456 503616
rect 446312 496868 446364 496874
rect 446312 496810 446364 496816
rect 446128 494624 446180 494630
rect 446128 494566 446180 494572
rect 445944 491292 445996 491298
rect 445944 491234 445996 491240
rect 445864 491150 446076 491178
rect 445944 491088 445996 491094
rect 445944 491030 445996 491036
rect 445852 485852 445904 485858
rect 445852 485794 445904 485800
rect 445864 417178 445892 485794
rect 445956 427553 445984 491030
rect 446048 437986 446076 491150
rect 446036 437980 446088 437986
rect 446036 437922 446088 437928
rect 446048 437510 446076 437922
rect 446036 437504 446088 437510
rect 446036 437446 446088 437452
rect 446140 434450 446168 494566
rect 446220 494012 446272 494018
rect 446220 493954 446272 493960
rect 446232 493406 446260 493954
rect 446220 493400 446272 493406
rect 446220 493342 446272 493348
rect 446128 434444 446180 434450
rect 446128 434386 446180 434392
rect 446140 433770 446168 434386
rect 446128 433764 446180 433770
rect 446128 433706 446180 433712
rect 446232 432954 446260 493342
rect 446324 441386 446352 496810
rect 446416 493338 446444 503610
rect 446404 493332 446456 493338
rect 446404 493274 446456 493280
rect 446508 487898 446536 523670
rect 446496 487892 446548 487898
rect 446496 487834 446548 487840
rect 446312 441380 446364 441386
rect 446312 441322 446364 441328
rect 446324 440434 446352 441322
rect 446312 440428 446364 440434
rect 446312 440370 446364 440376
rect 446220 432948 446272 432954
rect 446220 432890 446272 432896
rect 445942 427544 445998 427553
rect 445942 427479 445998 427488
rect 445956 422294 445984 427479
rect 445956 422266 446352 422294
rect 445852 417172 445904 417178
rect 445852 417114 445904 417120
rect 445668 358760 445720 358766
rect 445668 358702 445720 358708
rect 445680 357921 445708 358702
rect 445666 357912 445722 357921
rect 445666 357847 445722 357856
rect 445576 357400 445628 357406
rect 445576 357342 445628 357348
rect 445484 357332 445536 357338
rect 445484 357274 445536 357280
rect 445496 357241 445524 357274
rect 445482 357232 445538 357241
rect 445482 357167 445538 357176
rect 445588 356833 445616 357342
rect 445574 356824 445630 356833
rect 445574 356759 445630 356768
rect 445574 354104 445630 354113
rect 445574 354039 445576 354048
rect 445628 354039 445630 354048
rect 445576 354010 445628 354016
rect 445574 353016 445630 353025
rect 445574 352951 445630 352960
rect 445588 352646 445616 352951
rect 445576 352640 445628 352646
rect 445576 352582 445628 352588
rect 445576 352504 445628 352510
rect 445574 352472 445576 352481
rect 445628 352472 445630 352481
rect 445574 352407 445630 352416
rect 445576 351960 445628 351966
rect 445574 351928 445576 351937
rect 445628 351928 445630 351937
rect 445574 351863 445630 351872
rect 445482 350296 445538 350305
rect 445482 350231 445484 350240
rect 445536 350231 445538 350240
rect 445484 350202 445536 350208
rect 445482 345536 445538 345545
rect 445482 345471 445538 345480
rect 445496 344214 445524 345471
rect 445484 344208 445536 344214
rect 445484 344150 445536 344156
rect 445482 340640 445538 340649
rect 445482 340575 445484 340584
rect 445536 340575 445538 340584
rect 445484 340546 445536 340552
rect 445680 306374 445708 357847
rect 446128 353864 446180 353870
rect 446128 353806 446180 353812
rect 446036 352640 446088 352646
rect 446036 352582 446088 352588
rect 445944 349716 445996 349722
rect 445944 349658 445996 349664
rect 445956 349353 445984 349658
rect 445942 349344 445998 349353
rect 445942 349279 445998 349288
rect 445852 347744 445904 347750
rect 445852 347686 445904 347692
rect 445864 347177 445892 347686
rect 445850 347168 445906 347177
rect 445850 347103 445906 347112
rect 445758 346080 445814 346089
rect 445758 346015 445814 346024
rect 445588 306346 445708 306374
rect 445588 298042 445616 306346
rect 445668 298104 445720 298110
rect 445668 298046 445720 298052
rect 445576 298036 445628 298042
rect 445576 297978 445628 297984
rect 445392 297288 445444 297294
rect 445392 297230 445444 297236
rect 445404 296714 445432 297230
rect 445680 297022 445708 298046
rect 445668 297016 445720 297022
rect 445668 296958 445720 296964
rect 445404 296686 445616 296714
rect 445208 295996 445260 296002
rect 445208 295938 445260 295944
rect 445220 247926 445248 295938
rect 445392 295248 445444 295254
rect 445390 295216 445392 295225
rect 445444 295216 445446 295225
rect 445390 295151 445446 295160
rect 445484 295180 445536 295186
rect 445484 295122 445536 295128
rect 445496 294137 445524 295122
rect 445482 294128 445538 294137
rect 445482 294063 445538 294072
rect 445482 290592 445538 290601
rect 445482 290527 445538 290536
rect 445496 290426 445524 290527
rect 445484 290420 445536 290426
rect 445484 290362 445536 290368
rect 445484 280628 445536 280634
rect 445484 280570 445536 280576
rect 445496 280265 445524 280570
rect 445482 280256 445538 280265
rect 445482 280191 445538 280200
rect 445298 280120 445354 280129
rect 445298 280055 445354 280064
rect 445312 279041 445340 280055
rect 445298 279032 445354 279041
rect 445298 278967 445354 278976
rect 445208 247920 445260 247926
rect 445208 247862 445260 247868
rect 445208 240100 445260 240106
rect 445208 240042 445260 240048
rect 445220 239426 445248 240042
rect 445208 239420 445260 239426
rect 445208 239362 445260 239368
rect 445116 230444 445168 230450
rect 445116 230386 445168 230392
rect 445116 224256 445168 224262
rect 445116 224198 445168 224204
rect 445128 213353 445156 224198
rect 445114 213344 445170 213353
rect 445114 213279 445170 213288
rect 445128 212906 445156 213279
rect 445116 212900 445168 212906
rect 445116 212842 445168 212848
rect 445024 212424 445076 212430
rect 445024 212366 445076 212372
rect 445114 212392 445170 212401
rect 445114 212327 445116 212336
rect 445168 212327 445170 212336
rect 445116 212298 445168 212304
rect 445114 209536 445170 209545
rect 445114 209471 445170 209480
rect 445128 209098 445156 209471
rect 445116 209092 445168 209098
rect 445116 209034 445168 209040
rect 445114 208448 445170 208457
rect 445114 208383 445170 208392
rect 445128 208350 445156 208383
rect 445116 208344 445168 208350
rect 445116 208286 445168 208292
rect 445128 206938 445156 208286
rect 445036 206910 445156 206938
rect 444930 198792 444986 198801
rect 444930 198727 444986 198736
rect 444932 197804 444984 197810
rect 444932 197746 444984 197752
rect 444840 167680 444892 167686
rect 444840 167622 444892 167628
rect 444852 167346 444880 167622
rect 444840 167340 444892 167346
rect 444840 167282 444892 167288
rect 444656 163804 444708 163810
rect 444656 163746 444708 163752
rect 444668 163538 444696 163746
rect 444656 163532 444708 163538
rect 444656 163474 444708 163480
rect 444564 154556 444616 154562
rect 444564 154498 444616 154504
rect 444748 154556 444800 154562
rect 444748 154498 444800 154504
rect 444656 154420 444708 154426
rect 444656 154362 444708 154368
rect 444668 153678 444696 154362
rect 444760 153882 444788 154498
rect 444840 154352 444892 154358
rect 444840 154294 444892 154300
rect 444748 153876 444800 153882
rect 444748 153818 444800 153824
rect 444656 153672 444708 153678
rect 444656 153614 444708 153620
rect 444668 140865 444696 153614
rect 444852 153610 444880 154294
rect 444840 153604 444892 153610
rect 444840 153546 444892 153552
rect 444748 152040 444800 152046
rect 444748 151982 444800 151988
rect 444760 151706 444788 151982
rect 444748 151700 444800 151706
rect 444748 151642 444800 151648
rect 444852 144265 444880 153546
rect 444838 144256 444894 144265
rect 444838 144191 444894 144200
rect 444654 140856 444710 140865
rect 444654 140791 444710 140800
rect 444470 129840 444526 129849
rect 444470 129775 444526 129784
rect 444840 129056 444892 129062
rect 444840 128998 444892 129004
rect 443366 128752 443422 128761
rect 443366 128687 443422 128696
rect 443380 127634 443408 128687
rect 444852 128081 444880 128998
rect 444838 128072 444894 128081
rect 444838 128007 444894 128016
rect 444944 127634 444972 197746
rect 445036 169697 445064 206910
rect 445114 206816 445170 206825
rect 445114 206751 445170 206760
rect 445128 171086 445156 206751
rect 445220 201385 445248 239362
rect 445312 233918 445340 278967
rect 445390 275632 445446 275641
rect 445390 275567 445446 275576
rect 445300 233912 445352 233918
rect 445300 233854 445352 233860
rect 445206 201376 445262 201385
rect 445206 201311 445262 201320
rect 445312 201249 445340 233854
rect 445404 228410 445432 275567
rect 445484 269816 445536 269822
rect 445482 269784 445484 269793
rect 445536 269784 445538 269793
rect 445482 269719 445538 269728
rect 445482 268696 445538 268705
rect 445482 268631 445538 268640
rect 445496 268530 445524 268631
rect 445484 268524 445536 268530
rect 445484 268466 445536 268472
rect 445484 268388 445536 268394
rect 445484 268330 445536 268336
rect 445392 228404 445444 228410
rect 445392 228346 445444 228352
rect 445298 201240 445354 201249
rect 445298 201175 445354 201184
rect 445404 200122 445432 228346
rect 445208 200116 445260 200122
rect 445208 200058 445260 200064
rect 445392 200116 445444 200122
rect 445392 200058 445444 200064
rect 445220 198937 445248 200058
rect 445496 200002 445524 268330
rect 445588 224330 445616 296686
rect 445576 224324 445628 224330
rect 445576 224266 445628 224272
rect 445680 224262 445708 296958
rect 445772 281314 445800 346015
rect 445864 283665 445892 347103
rect 445956 288289 445984 349279
rect 446048 296546 446076 352582
rect 446140 297566 446168 353806
rect 446220 353388 446272 353394
rect 446220 353330 446272 353336
rect 446232 346662 446260 353330
rect 446324 347750 446352 422266
rect 446508 420986 446536 487834
rect 446600 486062 446628 561138
rect 447140 557660 447192 557666
rect 447140 557602 447192 557608
rect 447152 499574 447180 557602
rect 447796 512718 447824 583850
rect 447876 579692 447928 579698
rect 447876 579634 447928 579640
rect 447888 517886 447916 579634
rect 448152 578468 448204 578474
rect 448152 578410 448204 578416
rect 447968 574116 448020 574122
rect 447968 574058 448020 574064
rect 447876 517880 447928 517886
rect 447876 517822 447928 517828
rect 447980 514842 448008 574058
rect 448060 571532 448112 571538
rect 448060 571474 448112 571480
rect 448072 520946 448100 571474
rect 448164 541686 448192 578410
rect 448244 575544 448296 575550
rect 448244 575486 448296 575492
rect 448152 541680 448204 541686
rect 448152 541622 448204 541628
rect 448060 520940 448112 520946
rect 448060 520882 448112 520888
rect 447888 514826 448008 514842
rect 447876 514820 448008 514826
rect 447928 514814 448008 514820
rect 447876 514762 447928 514768
rect 447784 512712 447836 512718
rect 447784 512654 447836 512660
rect 447796 499574 447824 512654
rect 447888 503674 447916 514762
rect 447876 503668 447928 503674
rect 447876 503610 447928 503616
rect 447152 499546 447364 499574
rect 447140 496868 447192 496874
rect 447140 496810 447192 496816
rect 446956 493332 447008 493338
rect 446956 493274 447008 493280
rect 446588 486056 446640 486062
rect 446588 485998 446640 486004
rect 446600 485858 446628 485998
rect 446588 485852 446640 485858
rect 446588 485794 446640 485800
rect 446680 437504 446732 437510
rect 446680 437446 446732 437452
rect 446588 436756 446640 436762
rect 446588 436698 446640 436704
rect 446496 420980 446548 420986
rect 446496 420922 446548 420928
rect 446508 420646 446536 420922
rect 446496 420640 446548 420646
rect 446496 420582 446548 420588
rect 446496 417172 446548 417178
rect 446496 417114 446548 417120
rect 446508 380186 446536 417114
rect 446496 380180 446548 380186
rect 446496 380122 446548 380128
rect 446508 379574 446536 380122
rect 446496 379568 446548 379574
rect 446496 379510 446548 379516
rect 446600 373994 446628 436698
rect 446692 378146 446720 437446
rect 446864 433764 446916 433770
rect 446864 433706 446916 433712
rect 446772 432948 446824 432954
rect 446772 432890 446824 432896
rect 446784 381546 446812 432890
rect 446876 389230 446904 433706
rect 446968 431118 446996 493274
rect 447152 491230 447180 496810
rect 447140 491224 447192 491230
rect 447140 491166 447192 491172
rect 447336 485110 447364 499546
rect 447520 499546 447824 499574
rect 447520 497010 447548 499546
rect 447508 497004 447560 497010
rect 447508 496946 447560 496952
rect 447416 488776 447468 488782
rect 447416 488718 447468 488724
rect 447324 485104 447376 485110
rect 447324 485046 447376 485052
rect 447336 484634 447364 485046
rect 447324 484628 447376 484634
rect 447324 484570 447376 484576
rect 447140 439068 447192 439074
rect 447140 439010 447192 439016
rect 446956 431112 447008 431118
rect 446956 431054 447008 431060
rect 446864 389224 446916 389230
rect 446864 389166 446916 389172
rect 446772 381540 446824 381546
rect 446772 381482 446824 381488
rect 446680 378140 446732 378146
rect 446680 378082 446732 378088
rect 446508 373966 446628 373994
rect 446508 371278 446536 373966
rect 446496 371272 446548 371278
rect 446496 371214 446548 371220
rect 446508 351422 446536 371214
rect 446496 351416 446548 351422
rect 446496 351358 446548 351364
rect 446784 349722 446812 381482
rect 447048 379568 447100 379574
rect 447048 379510 447100 379516
rect 446772 349716 446824 349722
rect 446772 349658 446824 349664
rect 446312 347744 446364 347750
rect 446312 347686 446364 347692
rect 446404 346724 446456 346730
rect 446404 346666 446456 346672
rect 446220 346656 446272 346662
rect 446220 346598 446272 346604
rect 446232 313954 446260 346598
rect 446416 340882 446444 346666
rect 447060 342310 447088 379510
rect 447152 352510 447180 439010
rect 447336 413710 447364 484570
rect 447428 426902 447456 488718
rect 447520 440298 447548 496946
rect 448072 491094 448100 520882
rect 448164 494630 448192 541622
rect 448256 536110 448284 575486
rect 449164 568608 449216 568614
rect 449164 568550 449216 568556
rect 448244 536104 448296 536110
rect 448244 536046 448296 536052
rect 448152 494624 448204 494630
rect 448152 494566 448204 494572
rect 448256 494018 448284 536046
rect 449176 526454 449204 568550
rect 450544 563100 450596 563106
rect 450544 563042 450596 563048
rect 449256 555484 449308 555490
rect 449256 555426 449308 555432
rect 449164 526448 449216 526454
rect 449164 526390 449216 526396
rect 448428 517880 448480 517886
rect 448428 517822 448480 517828
rect 448440 517546 448468 517822
rect 448428 517540 448480 517546
rect 448428 517482 448480 517488
rect 448440 505102 448468 517482
rect 449164 507816 449216 507822
rect 449164 507758 449216 507764
rect 448520 505912 448572 505918
rect 448520 505854 448572 505860
rect 448428 505096 448480 505102
rect 448428 505038 448480 505044
rect 448244 494012 448296 494018
rect 448244 493954 448296 493960
rect 448060 491088 448112 491094
rect 448060 491030 448112 491036
rect 447692 484220 447744 484226
rect 447692 484162 447744 484168
rect 447508 440292 447560 440298
rect 447508 440234 447560 440240
rect 447416 426896 447468 426902
rect 447416 426838 447468 426844
rect 447600 414860 447652 414866
rect 447600 414802 447652 414808
rect 447324 413704 447376 413710
rect 447324 413646 447376 413652
rect 447336 412634 447364 413646
rect 447244 412606 447364 412634
rect 447140 352504 447192 352510
rect 447140 352446 447192 352452
rect 447048 342304 447100 342310
rect 447100 342252 447180 342258
rect 447048 342246 447180 342252
rect 447060 342230 447180 342246
rect 447060 342181 447088 342230
rect 446404 340876 446456 340882
rect 446404 340818 446456 340824
rect 446220 313948 446272 313954
rect 446220 313890 446272 313896
rect 446128 297560 446180 297566
rect 446128 297502 446180 297508
rect 446036 296540 446088 296546
rect 446036 296482 446088 296488
rect 445942 288280 445998 288289
rect 445942 288215 445998 288224
rect 445956 287502 445984 288215
rect 445944 287496 445996 287502
rect 445944 287438 445996 287444
rect 445850 283656 445906 283665
rect 445850 283591 445906 283600
rect 445864 282946 445892 283591
rect 445852 282940 445904 282946
rect 445852 282882 445904 282888
rect 446232 282878 446260 313890
rect 446416 284850 446444 340818
rect 446494 291816 446550 291825
rect 446494 291751 446550 291760
rect 446404 284844 446456 284850
rect 446404 284786 446456 284792
rect 446220 282872 446272 282878
rect 446220 282814 446272 282820
rect 445760 281308 445812 281314
rect 445760 281250 445812 281256
rect 445760 268524 445812 268530
rect 445760 268466 445812 268472
rect 445668 224256 445720 224262
rect 445668 224198 445720 224204
rect 445666 223000 445722 223009
rect 445666 222935 445722 222944
rect 445574 222456 445630 222465
rect 445574 222391 445630 222400
rect 445588 222290 445616 222391
rect 445576 222284 445628 222290
rect 445576 222226 445628 222232
rect 445680 222222 445708 222935
rect 445668 222216 445720 222222
rect 445668 222158 445720 222164
rect 445574 221368 445630 221377
rect 445574 221303 445630 221312
rect 445588 220862 445616 221303
rect 445576 220856 445628 220862
rect 445576 220798 445628 220804
rect 445666 220824 445722 220833
rect 445666 220759 445722 220768
rect 445574 219736 445630 219745
rect 445574 219671 445630 219680
rect 445588 219502 445616 219671
rect 445680 219638 445708 220759
rect 445668 219632 445720 219638
rect 445668 219574 445720 219580
rect 445576 219496 445628 219502
rect 445576 219438 445628 219444
rect 445772 209774 445800 268466
rect 446416 229770 446444 284786
rect 446508 243574 446536 291751
rect 446680 287496 446732 287502
rect 446680 287438 446732 287444
rect 446588 282940 446640 282946
rect 446588 282882 446640 282888
rect 446496 243568 446548 243574
rect 446496 243510 446548 243516
rect 446496 241460 446548 241466
rect 446496 241402 446548 241408
rect 446508 240786 446536 241402
rect 446496 240780 446548 240786
rect 446496 240722 446548 240728
rect 446404 229764 446456 229770
rect 446404 229706 446456 229712
rect 445944 225072 445996 225078
rect 445944 225014 445996 225020
rect 445852 225004 445904 225010
rect 445852 224946 445904 224952
rect 445864 216481 445892 224946
rect 445956 217326 445984 225014
rect 445944 217320 445996 217326
rect 445944 217262 445996 217268
rect 445956 217025 445984 217262
rect 445942 217016 445998 217025
rect 445942 216951 445998 216960
rect 445850 216472 445906 216481
rect 445850 216407 445906 216416
rect 445864 215966 445892 216407
rect 445852 215960 445904 215966
rect 445852 215902 445904 215908
rect 446036 215892 446088 215898
rect 446036 215834 446088 215840
rect 445944 212900 445996 212906
rect 445944 212842 445996 212848
rect 445772 209746 445892 209774
rect 445668 209160 445720 209166
rect 445668 209102 445720 209108
rect 445680 209001 445708 209102
rect 445666 208992 445722 209001
rect 445666 208927 445722 208936
rect 445666 207904 445722 207913
rect 445666 207839 445722 207848
rect 445680 207670 445708 207839
rect 445668 207664 445720 207670
rect 445668 207606 445720 207612
rect 445574 204232 445630 204241
rect 445574 204167 445630 204176
rect 445312 199974 445524 200002
rect 445206 198928 445262 198937
rect 445206 198863 445262 198872
rect 445312 198257 445340 199974
rect 445482 199880 445538 199889
rect 445482 199815 445538 199824
rect 445298 198248 445354 198257
rect 445298 198183 445354 198192
rect 445312 198082 445340 198183
rect 445300 198076 445352 198082
rect 445300 198018 445352 198024
rect 445312 197810 445340 198018
rect 445300 197804 445352 197810
rect 445300 197746 445352 197752
rect 445298 197704 445354 197713
rect 445298 197639 445354 197648
rect 445312 197402 445340 197639
rect 445300 197396 445352 197402
rect 445300 197338 445352 197344
rect 445392 197260 445444 197266
rect 445392 197202 445444 197208
rect 445208 197192 445260 197198
rect 445208 197134 445260 197140
rect 445116 171080 445168 171086
rect 445116 171022 445168 171028
rect 445022 169688 445078 169697
rect 445022 169623 445078 169632
rect 445116 168360 445168 168366
rect 445116 168302 445168 168308
rect 445024 167340 445076 167346
rect 445024 167282 445076 167288
rect 445036 135318 445064 167282
rect 445128 153746 445156 168302
rect 445220 162858 445248 197134
rect 445404 196625 445432 197202
rect 445496 197198 445524 199815
rect 445484 197192 445536 197198
rect 445484 197134 445536 197140
rect 445588 196654 445616 204167
rect 445666 202600 445722 202609
rect 445722 202558 445800 202586
rect 445666 202535 445722 202544
rect 445668 201544 445720 201550
rect 445666 201512 445668 201521
rect 445720 201512 445722 201521
rect 445666 201447 445722 201456
rect 445772 197334 445800 202558
rect 445760 197328 445812 197334
rect 445760 197270 445812 197276
rect 445666 197160 445722 197169
rect 445666 197095 445722 197104
rect 445576 196648 445628 196654
rect 445390 196616 445446 196625
rect 445576 196590 445628 196596
rect 445390 196551 445446 196560
rect 445680 196042 445708 197095
rect 445772 196110 445800 197270
rect 445864 196217 445892 209746
rect 445850 196208 445906 196217
rect 445850 196143 445906 196152
rect 445760 196104 445812 196110
rect 445760 196046 445812 196052
rect 445668 196036 445720 196042
rect 445668 195978 445720 195984
rect 445864 180794 445892 196143
rect 445956 195294 445984 212842
rect 445944 195288 445996 195294
rect 445944 195230 445996 195236
rect 446048 190454 446076 215834
rect 446416 203998 446444 229706
rect 446404 203992 446456 203998
rect 446404 203934 446456 203940
rect 446508 202774 446536 240722
rect 446600 236706 446628 282882
rect 446692 247722 446720 287438
rect 446772 281308 446824 281314
rect 446772 281250 446824 281256
rect 446680 247716 446732 247722
rect 446680 247658 446732 247664
rect 446588 236700 446640 236706
rect 446588 236642 446640 236648
rect 446600 203386 446628 236642
rect 446692 205358 446720 247658
rect 446784 241466 446812 281250
rect 447152 273222 447180 342230
rect 447244 340610 447272 412606
rect 447416 389224 447468 389230
rect 447416 389166 447468 389172
rect 447428 350266 447456 389166
rect 447508 378140 447560 378146
rect 447508 378082 447560 378088
rect 447520 376786 447548 378082
rect 447508 376780 447560 376786
rect 447508 376722 447560 376728
rect 447520 351966 447548 376722
rect 447508 351960 447560 351966
rect 447508 351902 447560 351908
rect 447416 350260 447468 350266
rect 447416 350202 447468 350208
rect 447324 344208 447376 344214
rect 447324 344150 447376 344156
rect 447232 340604 447284 340610
rect 447232 340546 447284 340552
rect 447140 273216 447192 273222
rect 447140 273158 447192 273164
rect 447244 269822 447272 340546
rect 447336 280634 447364 344150
rect 447428 290426 447456 350202
rect 447520 295186 447548 351902
rect 447612 342242 447640 414802
rect 447704 412622 447732 484162
rect 447876 440428 447928 440434
rect 447876 440370 447928 440376
rect 447784 440292 447836 440298
rect 447784 440234 447836 440240
rect 447692 412616 447744 412622
rect 447692 412558 447744 412564
rect 447704 412010 447732 412558
rect 447692 412004 447744 412010
rect 447692 411946 447744 411952
rect 447796 366994 447824 440234
rect 447888 369170 447916 440370
rect 447968 426896 448020 426902
rect 447968 426838 448020 426844
rect 447980 376038 448008 426838
rect 448532 384334 448560 505854
rect 448612 504416 448664 504422
rect 448612 504358 448664 504364
rect 448624 385694 448652 504358
rect 448796 491700 448848 491706
rect 448796 491642 448848 491648
rect 448808 487354 448836 491642
rect 448796 487348 448848 487354
rect 448796 487290 448848 487296
rect 448704 487212 448756 487218
rect 448704 487154 448756 487160
rect 448716 484362 448744 487154
rect 448704 484356 448756 484362
rect 448704 484298 448756 484304
rect 448808 470594 448836 487290
rect 448716 470566 448836 470594
rect 448716 419490 448744 470566
rect 448704 419484 448756 419490
rect 448704 419426 448756 419432
rect 449176 388482 449204 507758
rect 449268 505918 449296 555426
rect 449348 526448 449400 526454
rect 449348 526390 449400 526396
rect 449256 505912 449308 505918
rect 449256 505854 449308 505860
rect 449256 497820 449308 497826
rect 449256 497762 449308 497768
rect 449268 412622 449296 497762
rect 449360 496874 449388 526390
rect 450556 522374 450584 563042
rect 454684 556912 454736 556918
rect 454684 556854 454736 556860
rect 450544 522368 450596 522374
rect 450544 522310 450596 522316
rect 450556 518894 450584 522310
rect 454696 522306 454724 556854
rect 456708 555552 456760 555558
rect 456708 555494 456760 555500
rect 454040 522300 454092 522306
rect 454040 522242 454092 522248
rect 454684 522300 454736 522306
rect 454684 522242 454736 522248
rect 450556 518866 450676 518894
rect 450176 508564 450228 508570
rect 450176 508506 450228 508512
rect 450084 507204 450136 507210
rect 450084 507146 450136 507152
rect 449992 507136 450044 507142
rect 449992 507078 450044 507084
rect 449900 505164 449952 505170
rect 449900 505106 449952 505112
rect 449912 505034 449940 505106
rect 449900 505028 449952 505034
rect 449900 504970 449952 504976
rect 450004 504506 450032 507078
rect 449912 504478 450032 504506
rect 449348 496868 449400 496874
rect 449348 496810 449400 496816
rect 449348 484356 449400 484362
rect 449348 484298 449400 484304
rect 449360 420918 449388 484298
rect 449440 420980 449492 420986
rect 449440 420922 449492 420928
rect 449348 420912 449400 420918
rect 449348 420854 449400 420860
rect 449256 412616 449308 412622
rect 449256 412558 449308 412564
rect 448704 388476 448756 388482
rect 448704 388418 448756 388424
rect 449164 388476 449216 388482
rect 449164 388418 449216 388424
rect 448612 385688 448664 385694
rect 448612 385630 448664 385636
rect 448520 384328 448572 384334
rect 448520 384270 448572 384276
rect 447968 376032 448020 376038
rect 447968 375974 448020 375980
rect 447876 369164 447928 369170
rect 447876 369106 447928 369112
rect 447784 366988 447836 366994
rect 447784 366930 447836 366936
rect 447888 353870 447916 369106
rect 447876 353864 447928 353870
rect 447876 353806 447928 353812
rect 447980 353394 448008 375974
rect 448532 361554 448560 384270
rect 448520 361548 448572 361554
rect 448520 361490 448572 361496
rect 448624 360194 448652 385630
rect 448716 365702 448744 388418
rect 448704 365696 448756 365702
rect 448704 365638 448756 365644
rect 448612 360188 448664 360194
rect 448612 360130 448664 360136
rect 449268 354074 449296 412558
rect 449452 373994 449480 420922
rect 449360 373966 449480 373994
rect 449360 373318 449388 373966
rect 449348 373312 449400 373318
rect 449348 373254 449400 373260
rect 448428 354068 448480 354074
rect 448428 354010 448480 354016
rect 449256 354068 449308 354074
rect 449256 354010 449308 354016
rect 447968 353388 448020 353394
rect 447968 353330 448020 353336
rect 447600 342236 447652 342242
rect 447600 342178 447652 342184
rect 447612 340950 447640 342178
rect 447600 340944 447652 340950
rect 447600 340886 447652 340892
rect 448440 297362 448468 354010
rect 449164 353320 449216 353326
rect 449164 353262 449216 353268
rect 448612 352504 448664 352510
rect 448612 352446 448664 352452
rect 448428 297356 448480 297362
rect 448428 297298 448480 297304
rect 448440 296714 448468 297298
rect 448440 296686 448560 296714
rect 447508 295180 447560 295186
rect 447508 295122 447560 295128
rect 447520 294642 447548 295122
rect 447508 294636 447560 294642
rect 447508 294578 447560 294584
rect 447416 290420 447468 290426
rect 447416 290362 447468 290368
rect 447968 290420 448020 290426
rect 447968 290362 448020 290368
rect 447876 289876 447928 289882
rect 447876 289818 447928 289824
rect 447784 287156 447836 287162
rect 447784 287098 447836 287104
rect 447324 280628 447376 280634
rect 447324 280570 447376 280576
rect 447232 269816 447284 269822
rect 447232 269758 447284 269764
rect 447244 258074 447272 269758
rect 447152 258046 447272 258074
rect 446864 243568 446916 243574
rect 446864 243510 446916 243516
rect 446772 241460 446824 241466
rect 446772 241402 446824 241408
rect 446876 206825 446904 243510
rect 446862 206816 446918 206825
rect 446862 206751 446918 206760
rect 446680 205352 446732 205358
rect 446680 205294 446732 205300
rect 446588 203380 446640 203386
rect 446588 203322 446640 203328
rect 446496 202768 446548 202774
rect 446496 202710 446548 202716
rect 447152 197266 447180 258046
rect 447796 226370 447824 287098
rect 447888 233238 447916 289818
rect 447980 235278 448008 290362
rect 448060 280628 448112 280634
rect 448060 280570 448112 280576
rect 447968 235272 448020 235278
rect 447968 235214 448020 235220
rect 447876 233232 447928 233238
rect 447876 233174 447928 233180
rect 447876 227792 447928 227798
rect 447876 227734 447928 227740
rect 447784 226364 447836 226370
rect 447784 226306 447836 226312
rect 447796 204814 447824 226306
rect 447784 204808 447836 204814
rect 447784 204750 447836 204756
rect 447888 202842 447916 227734
rect 447980 205630 448008 235214
rect 448072 228478 448100 280570
rect 448152 233232 448204 233238
rect 448152 233174 448204 233180
rect 448164 231878 448192 233174
rect 448152 231872 448204 231878
rect 448152 231814 448204 231820
rect 448060 228472 448112 228478
rect 448060 228414 448112 228420
rect 448072 227798 448100 228414
rect 448060 227792 448112 227798
rect 448060 227734 448112 227740
rect 448164 205902 448192 231814
rect 448532 211138 448560 296686
rect 448624 295254 448652 352446
rect 448612 295248 448664 295254
rect 448612 295190 448664 295196
rect 448624 294030 448652 295190
rect 448612 294024 448664 294030
rect 448612 293966 448664 293972
rect 449176 267714 449204 353262
rect 449360 343942 449388 373254
rect 449912 369918 449940 504478
rect 450096 504370 450124 507146
rect 450004 504342 450124 504370
rect 450004 395350 450032 504342
rect 450188 489914 450216 508506
rect 450544 505028 450596 505034
rect 450544 504970 450596 504976
rect 450096 489886 450216 489914
rect 450096 398138 450124 489886
rect 450084 398132 450136 398138
rect 450084 398074 450136 398080
rect 449992 395344 450044 395350
rect 449992 395286 450044 395292
rect 449900 369912 449952 369918
rect 449900 369854 449952 369860
rect 450004 363866 450032 395286
rect 450096 364342 450124 398074
rect 450556 393990 450584 504970
rect 450648 491706 450676 518866
rect 452660 509992 452712 509998
rect 452660 509934 452712 509940
rect 451280 509924 451332 509930
rect 451280 509866 451332 509872
rect 450636 491700 450688 491706
rect 450636 491642 450688 491648
rect 450544 393984 450596 393990
rect 450544 393926 450596 393932
rect 450556 393314 450584 393926
rect 450188 393286 450584 393314
rect 450084 364336 450136 364342
rect 450084 364278 450136 364284
rect 449992 363860 450044 363866
rect 449992 363802 450044 363808
rect 450188 362914 450216 393286
rect 451292 364410 451320 509866
rect 452672 365770 452700 509934
rect 452752 505096 452804 505102
rect 452752 505038 452804 505044
rect 452764 494086 452792 505038
rect 454052 499526 454080 522242
rect 456720 500818 456748 555494
rect 458180 504484 458232 504490
rect 458180 504426 458232 504432
rect 458192 503742 458220 504426
rect 458180 503736 458232 503742
rect 458180 503678 458232 503684
rect 458824 503736 458876 503742
rect 458824 503678 458876 503684
rect 456708 500812 456760 500818
rect 456708 500754 456760 500760
rect 456720 500410 456748 500754
rect 456708 500404 456760 500410
rect 456708 500346 456760 500352
rect 457444 500404 457496 500410
rect 457444 500346 457496 500352
rect 454040 499520 454092 499526
rect 454040 499462 454092 499468
rect 452752 494080 452804 494086
rect 452752 494022 452804 494028
rect 457456 441862 457484 500346
rect 458836 442338 458864 503678
rect 459560 501628 459612 501634
rect 459560 501570 459612 501576
rect 460204 501628 460256 501634
rect 460204 501570 460256 501576
rect 459572 501022 459600 501570
rect 459560 501016 459612 501022
rect 459560 500958 459612 500964
rect 458824 442332 458876 442338
rect 458824 442274 458876 442280
rect 460216 442270 460244 501570
rect 460204 442264 460256 442270
rect 460204 442206 460256 442212
rect 457444 441856 457496 441862
rect 457444 441798 457496 441804
rect 455328 367940 455380 367946
rect 455328 367882 455380 367888
rect 455340 366994 455368 367882
rect 454040 366988 454092 366994
rect 454040 366930 454092 366936
rect 455328 366988 455380 366994
rect 455328 366930 455380 366936
rect 452660 365764 452712 365770
rect 452660 365706 452712 365712
rect 451280 364404 451332 364410
rect 451280 364346 451332 364352
rect 450176 362908 450228 362914
rect 450176 362850 450228 362856
rect 454052 352646 454080 366930
rect 457456 355366 457484 441798
rect 458824 411936 458876 411942
rect 458824 411878 458876 411884
rect 458836 357338 458864 411878
rect 458824 357332 458876 357338
rect 458824 357274 458876 357280
rect 457444 355360 457496 355366
rect 457444 355302 457496 355308
rect 454040 352640 454092 352646
rect 454040 352582 454092 352588
rect 449348 343936 449400 343942
rect 449348 343878 449400 343884
rect 461596 307154 461624 699654
rect 489184 584520 489236 584526
rect 489184 584462 489236 584468
rect 485044 584452 485096 584458
rect 485044 584394 485096 584400
rect 483664 584112 483716 584118
rect 483664 584054 483716 584060
rect 482284 555688 482336 555694
rect 482284 555630 482336 555636
rect 464344 555620 464396 555626
rect 464344 555562 464396 555568
rect 464356 504490 464384 555562
rect 464344 504484 464396 504490
rect 464344 504426 464396 504432
rect 482296 500886 482324 555630
rect 483676 512786 483704 584054
rect 483664 512780 483716 512786
rect 483664 512722 483716 512728
rect 485056 511970 485084 584394
rect 486424 556980 486476 556986
rect 486424 556922 486476 556928
rect 485044 511964 485096 511970
rect 485044 511906 485096 511912
rect 486436 501634 486464 556922
rect 489196 509998 489224 584462
rect 493324 584248 493376 584254
rect 493324 584190 493376 584196
rect 490564 584180 490616 584186
rect 490564 584122 490616 584128
rect 489184 509992 489236 509998
rect 489184 509934 489236 509940
rect 490576 509930 490604 584122
rect 490564 509924 490616 509930
rect 490564 509866 490616 509872
rect 493336 508570 493364 584190
rect 493324 508564 493376 508570
rect 493324 508506 493376 508512
rect 486424 501628 486476 501634
rect 486424 501570 486476 501576
rect 482284 500880 482336 500886
rect 482284 500822 482336 500828
rect 466828 498840 466880 498846
rect 466828 498782 466880 498788
rect 467748 498840 467800 498846
rect 467748 498782 467800 498788
rect 466840 498234 466868 498782
rect 466828 498228 466880 498234
rect 466828 498170 466880 498176
rect 467760 442950 467788 498782
rect 467104 442944 467156 442950
rect 467104 442886 467156 442892
rect 467748 442944 467800 442950
rect 467748 442886 467800 442892
rect 467116 441930 467144 442886
rect 467104 441924 467156 441930
rect 467104 441866 467156 441872
rect 467116 354657 467144 441866
rect 472716 412004 472768 412010
rect 472716 411946 472768 411952
rect 472728 411330 472756 411946
rect 472716 411324 472768 411330
rect 472716 411266 472768 411272
rect 472728 393314 472756 411266
rect 472636 393286 472756 393314
rect 467102 354648 467158 354657
rect 467102 354583 467158 354592
rect 472636 340814 472664 393286
rect 472624 340808 472676 340814
rect 472624 340750 472676 340756
rect 472636 339522 472664 340750
rect 471244 339516 471296 339522
rect 471244 339458 471296 339464
rect 472624 339516 472676 339522
rect 472624 339458 472676 339464
rect 461584 307148 461636 307154
rect 461584 307090 461636 307096
rect 456064 294636 456116 294642
rect 456064 294578 456116 294584
rect 449256 294024 449308 294030
rect 449256 293966 449308 293972
rect 449164 267708 449216 267714
rect 449164 267650 449216 267656
rect 448520 211132 448572 211138
rect 448520 211074 448572 211080
rect 449176 211070 449204 267650
rect 449268 233306 449296 293966
rect 449348 268388 449400 268394
rect 449348 268330 449400 268336
rect 449360 267753 449388 268330
rect 449346 267744 449402 267753
rect 449346 267679 449402 267688
rect 449256 233300 449308 233306
rect 449256 233242 449308 233248
rect 449164 211064 449216 211070
rect 449164 211006 449216 211012
rect 449268 208350 449296 233242
rect 456076 225010 456104 294578
rect 471256 269074 471284 339458
rect 494072 304774 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 699718 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 526444 699712 526496 699718
rect 526444 699654 526496 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 513378 585440 513434 585449
rect 513378 585375 513434 585384
rect 513562 585440 513618 585449
rect 513562 585375 513564 585384
rect 513392 585342 513420 585375
rect 513616 585375 513618 585384
rect 513564 585346 513616 585352
rect 513380 585336 513432 585342
rect 513380 585278 513432 585284
rect 516416 585268 516468 585274
rect 516416 585210 516468 585216
rect 516138 584624 516194 584633
rect 516138 584559 516194 584568
rect 513932 584520 513984 584526
rect 513932 584462 513984 584468
rect 513564 584452 513616 584458
rect 513564 584394 513616 584400
rect 500224 584316 500276 584322
rect 500224 584258 500276 584264
rect 497464 583908 497516 583914
rect 497464 583850 497516 583856
rect 497476 507210 497504 583850
rect 497464 507204 497516 507210
rect 497464 507146 497516 507152
rect 500236 507142 500264 584258
rect 513380 584112 513432 584118
rect 513380 584054 513432 584060
rect 513288 583976 513340 583982
rect 513392 583953 513420 584054
rect 513576 583953 513604 584394
rect 513748 584384 513800 584390
rect 513748 584326 513800 584332
rect 513656 584180 513708 584186
rect 513656 584122 513708 584128
rect 513288 583918 513340 583924
rect 513378 583944 513434 583953
rect 513300 580145 513328 583918
rect 513562 583944 513618 583953
rect 513378 583879 513434 583888
rect 513472 583908 513524 583914
rect 513562 583879 513618 583888
rect 513472 583850 513524 583856
rect 513378 580544 513434 580553
rect 513378 580479 513434 580488
rect 513286 580136 513342 580145
rect 513286 580071 513342 580080
rect 502984 557116 503036 557122
rect 502984 557058 503036 557064
rect 501604 557048 501656 557054
rect 501604 556990 501656 556996
rect 500224 507136 500276 507142
rect 500224 507078 500276 507084
rect 501616 504422 501644 556990
rect 501604 504416 501656 504422
rect 501604 504358 501656 504364
rect 502996 498846 503024 557058
rect 513392 557002 513420 580479
rect 513484 579601 513512 583850
rect 513668 581777 513696 584122
rect 513760 582865 513788 584326
rect 513840 584248 513892 584254
rect 513840 584190 513892 584196
rect 513746 582856 513802 582865
rect 513746 582791 513802 582800
rect 513654 581768 513710 581777
rect 513654 581703 513710 581712
rect 513852 580689 513880 584190
rect 513944 582321 513972 584462
rect 516152 583778 516180 584559
rect 516324 584316 516376 584322
rect 516324 584258 516376 584264
rect 516232 584044 516284 584050
rect 516232 583986 516284 583992
rect 516140 583772 516192 583778
rect 516140 583714 516192 583720
rect 514850 582992 514906 583001
rect 514850 582927 514906 582936
rect 513930 582312 513986 582321
rect 513930 582247 513986 582256
rect 513838 580680 513894 580689
rect 513838 580615 513894 580624
rect 513470 579592 513526 579601
rect 513470 579527 513526 579536
rect 513470 577824 513526 577833
rect 513470 577759 513526 577768
rect 513484 557534 513512 577759
rect 513654 574152 513710 574161
rect 513654 574087 513710 574096
rect 513484 557506 513604 557534
rect 513392 556974 513512 557002
rect 513380 556844 513432 556850
rect 513380 556786 513432 556792
rect 513392 556481 513420 556786
rect 513378 556472 513434 556481
rect 513378 556407 513434 556416
rect 503732 556022 504942 556050
rect 503352 555960 503404 555966
rect 503352 555902 503404 555908
rect 503260 555892 503312 555898
rect 503260 555834 503312 555840
rect 503168 555824 503220 555830
rect 503168 555766 503220 555772
rect 503076 555756 503128 555762
rect 503076 555698 503128 555704
rect 503088 500954 503116 555698
rect 503180 502314 503208 555766
rect 503272 505102 503300 555834
rect 503364 507822 503392 555902
rect 503352 507816 503404 507822
rect 503352 507758 503404 507764
rect 503260 505096 503312 505102
rect 503260 505038 503312 505044
rect 503168 502308 503220 502314
rect 503168 502250 503220 502256
rect 503076 500948 503128 500954
rect 503076 500890 503128 500896
rect 503732 499574 503760 556022
rect 506860 554742 506888 556036
rect 507872 556022 508898 556050
rect 506848 554736 506900 554742
rect 506848 554678 506900 554684
rect 507872 514078 507900 556022
rect 510908 554130 510936 556036
rect 510896 554124 510948 554130
rect 510896 554066 510948 554072
rect 512932 553450 512960 556036
rect 513484 555966 513512 556974
rect 513472 555960 513524 555966
rect 513472 555902 513524 555908
rect 513576 555898 513604 557506
rect 513564 555892 513616 555898
rect 513564 555834 513616 555840
rect 513668 555830 513696 574087
rect 513746 573608 513802 573617
rect 513746 573543 513802 573552
rect 513656 555824 513708 555830
rect 513656 555766 513708 555772
rect 513760 555762 513788 573543
rect 513930 573064 513986 573073
rect 513930 572999 513986 573008
rect 513838 571432 513894 571441
rect 513838 571367 513894 571376
rect 513748 555756 513800 555762
rect 513748 555698 513800 555704
rect 513852 555558 513880 571367
rect 513944 556073 513972 572999
rect 513930 556064 513986 556073
rect 513930 555999 513986 556008
rect 513840 555552 513892 555558
rect 513840 555494 513892 555500
rect 512920 553444 512972 553450
rect 512920 553386 512972 553392
rect 514760 553444 514812 553450
rect 514760 553386 514812 553392
rect 507860 514072 507912 514078
rect 507860 514014 507912 514020
rect 513380 514072 513432 514078
rect 513380 514014 513432 514020
rect 513392 499574 513420 514014
rect 513748 512712 513800 512718
rect 513746 512680 513748 512689
rect 513800 512680 513802 512689
rect 513746 512615 513802 512624
rect 503732 499546 504496 499574
rect 513392 499546 513604 499574
rect 502984 498840 503036 498846
rect 502984 498782 503036 498788
rect 504468 484106 504496 499546
rect 513470 488744 513526 488753
rect 513470 488679 513526 488688
rect 513378 487520 513434 487529
rect 513378 487455 513434 487464
rect 513392 485790 513420 487455
rect 513484 486062 513512 488679
rect 513472 486056 513524 486062
rect 513472 485998 513524 486004
rect 513380 485784 513432 485790
rect 513380 485726 513432 485732
rect 513104 484288 513156 484294
rect 512946 484236 513104 484242
rect 512946 484230 513156 484236
rect 512946 484228 513144 484230
rect 512932 484214 513144 484228
rect 504468 484092 504942 484106
rect 504468 484078 504956 484092
rect 504928 482798 504956 484078
rect 506860 483002 506888 484092
rect 506848 482996 506900 483002
rect 506848 482938 506900 482944
rect 508884 482934 508912 484092
rect 508872 482928 508924 482934
rect 508872 482870 508924 482876
rect 504916 482792 504968 482798
rect 504916 482734 504968 482740
rect 510908 482322 510936 484092
rect 512932 482866 512960 484214
rect 513576 482934 513604 499546
rect 513746 485208 513802 485217
rect 513746 485143 513802 485152
rect 513760 485110 513788 485143
rect 513748 485104 513800 485110
rect 513748 485046 513800 485052
rect 514772 484294 514800 553386
rect 514864 512650 514892 582927
rect 516244 577017 516272 583986
rect 516336 578649 516364 584258
rect 516322 578640 516378 578649
rect 516322 578575 516378 578584
rect 516230 577008 516286 577017
rect 516230 576943 516286 576952
rect 516428 575521 516456 585210
rect 524420 583772 524472 583778
rect 524420 583714 524472 583720
rect 516690 577552 516746 577561
rect 516690 577487 516746 577496
rect 516414 575512 516470 575521
rect 516414 575447 516470 575456
rect 516506 572248 516562 572257
rect 516506 572183 516562 572192
rect 516322 571160 516378 571169
rect 516322 571095 516378 571104
rect 516230 569528 516286 569537
rect 516230 569463 516286 569472
rect 516138 568984 516194 568993
rect 516138 568919 516140 568928
rect 516192 568919 516194 568928
rect 516140 568890 516192 568896
rect 516244 568614 516272 569463
rect 516232 568608 516284 568614
rect 516232 568550 516284 568556
rect 516336 568426 516364 571095
rect 516414 570616 516470 570625
rect 516414 570551 516470 570560
rect 516152 568398 516364 568426
rect 516152 567474 516180 568398
rect 516428 568290 516456 570551
rect 516336 568262 516456 568290
rect 516230 567896 516286 567905
rect 516230 567831 516286 567840
rect 516060 567446 516180 567474
rect 516060 567202 516088 567446
rect 516244 567390 516272 567831
rect 516232 567384 516284 567390
rect 516138 567352 516194 567361
rect 516232 567326 516284 567332
rect 516138 567287 516140 567296
rect 516192 567287 516194 567296
rect 516140 567258 516192 567264
rect 516232 567248 516284 567254
rect 516060 567174 516180 567202
rect 516232 567190 516284 567196
rect 516152 557122 516180 567174
rect 516244 557534 516272 567190
rect 516336 564346 516364 568262
rect 516520 568154 516548 572183
rect 516598 570072 516654 570081
rect 516598 570007 516654 570016
rect 516428 568126 516548 568154
rect 516428 566930 516456 568126
rect 516508 568064 516560 568070
rect 516508 568006 516560 568012
rect 516520 567050 516548 568006
rect 516612 567186 516640 570007
rect 516600 567180 516652 567186
rect 516600 567122 516652 567128
rect 516508 567044 516560 567050
rect 516508 566986 516560 566992
rect 516428 566902 516640 566930
rect 516506 566808 516562 566817
rect 516506 566743 516562 566752
rect 516414 566264 516470 566273
rect 516414 566199 516470 566208
rect 516428 565894 516456 566199
rect 516520 566098 516548 566743
rect 516508 566092 516560 566098
rect 516508 566034 516560 566040
rect 516416 565888 516468 565894
rect 516416 565830 516468 565836
rect 516506 565312 516562 565321
rect 516506 565247 516562 565256
rect 516414 564768 516470 564777
rect 516520 564738 516548 565247
rect 516414 564703 516470 564712
rect 516508 564732 516560 564738
rect 516428 564534 516456 564703
rect 516508 564674 516560 564680
rect 516416 564528 516468 564534
rect 516416 564470 516468 564476
rect 516336 564318 516456 564346
rect 516322 564224 516378 564233
rect 516322 564159 516378 564168
rect 516336 563786 516364 564159
rect 516324 563780 516376 563786
rect 516324 563722 516376 563728
rect 516322 563680 516378 563689
rect 516322 563615 516378 563624
rect 516336 563310 516364 563615
rect 516324 563304 516376 563310
rect 516324 563246 516376 563252
rect 516322 563136 516378 563145
rect 516322 563071 516324 563080
rect 516376 563071 516378 563080
rect 516324 563042 516376 563048
rect 516322 562592 516378 562601
rect 516322 562527 516324 562536
rect 516376 562527 516378 562536
rect 516324 562498 516376 562504
rect 516322 562048 516378 562057
rect 516322 561983 516324 561992
rect 516376 561983 516378 561992
rect 516324 561954 516376 561960
rect 516322 561504 516378 561513
rect 516322 561439 516324 561448
rect 516376 561439 516378 561448
rect 516324 561410 516376 561416
rect 516322 559328 516378 559337
rect 516322 559263 516378 559272
rect 516336 559026 516364 559263
rect 516324 559020 516376 559026
rect 516324 558962 516376 558968
rect 516324 557728 516376 557734
rect 516322 557696 516324 557705
rect 516376 557696 516378 557705
rect 516322 557631 516378 557640
rect 516244 557506 516364 557534
rect 516230 557152 516286 557161
rect 516140 557116 516192 557122
rect 516230 557087 516286 557096
rect 516140 557058 516192 557064
rect 516138 556608 516194 556617
rect 516138 556543 516194 556552
rect 516152 556306 516180 556543
rect 516140 556300 516192 556306
rect 516140 556242 516192 556248
rect 516244 556238 516272 557087
rect 516336 557054 516364 557506
rect 516324 557048 516376 557054
rect 516324 556990 516376 556996
rect 516428 556918 516456 564318
rect 516506 559872 516562 559881
rect 516506 559807 516562 559816
rect 516520 558958 516548 559807
rect 516508 558952 516560 558958
rect 516508 558894 516560 558900
rect 516506 558784 516562 558793
rect 516506 558719 516562 558728
rect 516520 557802 516548 558719
rect 516508 557796 516560 557802
rect 516508 557738 516560 557744
rect 516612 557682 516640 566902
rect 516520 557654 516640 557682
rect 516416 556912 516468 556918
rect 516416 556854 516468 556860
rect 516232 556232 516284 556238
rect 516232 556174 516284 556180
rect 516520 555694 516548 557654
rect 516600 557592 516652 557598
rect 516600 557534 516652 557540
rect 516612 556986 516640 557534
rect 516600 556980 516652 556986
rect 516600 556922 516652 556928
rect 516508 555688 516560 555694
rect 516508 555630 516560 555636
rect 516704 555490 516732 577487
rect 516874 576464 516930 576473
rect 516874 576399 516930 576408
rect 516782 573336 516838 573345
rect 516782 573271 516838 573280
rect 516796 568070 516824 573271
rect 516784 568064 516836 568070
rect 516784 568006 516836 568012
rect 516888 567254 516916 576399
rect 516966 576056 517022 576065
rect 516966 575991 517022 576000
rect 516876 567248 516928 567254
rect 516876 567190 516928 567196
rect 516876 567112 516928 567118
rect 516876 567054 516928 567060
rect 516784 567044 516836 567050
rect 516784 566986 516836 566992
rect 516796 557666 516824 566986
rect 516784 557660 516836 557666
rect 516784 557602 516836 557608
rect 516888 556170 516916 567054
rect 516876 556164 516928 556170
rect 516876 556106 516928 556112
rect 516980 555626 517008 575991
rect 517426 574968 517482 574977
rect 517482 574926 517560 574954
rect 517426 574903 517482 574912
rect 517426 560960 517482 560969
rect 517426 560895 517482 560904
rect 517242 560416 517298 560425
rect 517242 560351 517298 560360
rect 517058 558240 517114 558249
rect 517058 558175 517114 558184
rect 517072 557666 517100 558175
rect 517060 557660 517112 557666
rect 517060 557602 517112 557608
rect 516968 555620 517020 555626
rect 516968 555562 517020 555568
rect 516692 555484 516744 555490
rect 516692 555426 516744 555432
rect 516784 554804 516836 554810
rect 516784 554746 516836 554752
rect 516416 517540 516468 517546
rect 516416 517482 516468 517488
rect 516140 516112 516192 516118
rect 516140 516054 516192 516060
rect 516152 514826 516180 516054
rect 516140 514820 516192 514826
rect 516140 514762 516192 514768
rect 516152 513346 516180 514762
rect 516152 513318 516364 513346
rect 516140 512780 516192 512786
rect 516140 512722 516192 512728
rect 514852 512644 514904 512650
rect 514852 512586 514904 512592
rect 516152 512417 516180 512722
rect 516138 512408 516194 512417
rect 516138 512343 516194 512352
rect 516138 510096 516194 510105
rect 516138 510031 516194 510040
rect 516152 509930 516180 510031
rect 516140 509924 516192 509930
rect 516140 509866 516192 509872
rect 516138 508872 516194 508881
rect 516138 508807 516140 508816
rect 516192 508807 516194 508816
rect 516140 508778 516192 508784
rect 516140 507816 516192 507822
rect 516140 507758 516192 507764
rect 516152 506569 516180 507758
rect 516138 506560 516194 506569
rect 516138 506495 516194 506504
rect 516140 505096 516192 505102
rect 516140 505038 516192 505044
rect 516152 504257 516180 505038
rect 516138 504248 516194 504257
rect 516138 504183 516194 504192
rect 516336 503169 516364 513318
rect 516428 507793 516456 517482
rect 516414 507784 516470 507793
rect 516414 507719 516470 507728
rect 516322 503160 516378 503169
rect 516322 503095 516378 503104
rect 516138 500848 516194 500857
rect 516138 500783 516140 500792
rect 516192 500783 516194 500792
rect 516140 500754 516192 500760
rect 516140 500540 516192 500546
rect 516140 500482 516192 500488
rect 516152 499633 516180 500482
rect 516138 499624 516194 499633
rect 516138 499559 516194 499568
rect 516138 498536 516194 498545
rect 516138 498471 516140 498480
rect 516192 498471 516194 498480
rect 516140 498442 516192 498448
rect 516140 498160 516192 498166
rect 516140 498102 516192 498108
rect 516152 497321 516180 498102
rect 516138 497312 516194 497321
rect 516138 497247 516194 497256
rect 516230 496224 516286 496233
rect 516230 496159 516286 496168
rect 516244 495514 516272 496159
rect 516232 495508 516284 495514
rect 516232 495450 516284 495456
rect 516232 494012 516284 494018
rect 516232 493954 516284 493960
rect 516244 492697 516272 493954
rect 516322 493912 516378 493921
rect 516322 493847 516378 493856
rect 516230 492688 516286 492697
rect 516140 492652 516192 492658
rect 516230 492623 516286 492632
rect 516140 492594 516192 492600
rect 516152 491609 516180 492594
rect 516138 491600 516194 491609
rect 516138 491535 516194 491544
rect 516140 491224 516192 491230
rect 516140 491166 516192 491172
rect 516152 490385 516180 491166
rect 516138 490376 516194 490385
rect 516138 490311 516194 490320
rect 516336 489914 516364 493847
rect 516244 489886 516364 489914
rect 516138 486976 516194 486985
rect 516138 486911 516194 486920
rect 516152 486470 516180 486911
rect 516140 486464 516192 486470
rect 516140 486406 516192 486412
rect 516140 485784 516192 485790
rect 516138 485752 516140 485761
rect 516192 485752 516194 485761
rect 516138 485687 516194 485696
rect 516244 484362 516272 489886
rect 516692 489864 516744 489870
rect 516692 489806 516744 489812
rect 516704 489297 516732 489806
rect 516690 489288 516746 489297
rect 516690 489223 516746 489232
rect 516232 484356 516284 484362
rect 516232 484298 516284 484304
rect 514760 484288 514812 484294
rect 514760 484230 514812 484236
rect 513564 482928 513616 482934
rect 513564 482870 513616 482876
rect 512920 482860 512972 482866
rect 512920 482802 512972 482808
rect 510896 482316 510948 482322
rect 510896 482258 510948 482264
rect 516796 460934 516824 554746
rect 517152 514072 517204 514078
rect 517152 514014 517204 514020
rect 517164 513505 517192 514014
rect 517150 513496 517206 513505
rect 517150 513431 517206 513440
rect 516966 505472 517022 505481
rect 516966 505407 516968 505416
rect 517020 505407 517022 505416
rect 516968 505378 517020 505384
rect 516874 501936 516930 501945
rect 516874 501871 516930 501880
rect 516888 501430 516916 501871
rect 516876 501424 516928 501430
rect 516876 501366 516928 501372
rect 516874 495000 516930 495009
rect 516874 494935 516930 494944
rect 516428 460906 516824 460934
rect 516428 460222 516456 460906
rect 516416 460216 516468 460222
rect 516416 460158 516468 460164
rect 513472 442332 513524 442338
rect 513472 442274 513524 442280
rect 513380 441788 513432 441794
rect 513380 441730 513432 441736
rect 513392 430681 513420 441730
rect 513484 432313 513512 442274
rect 516232 441652 516284 441658
rect 516284 441600 516364 441614
rect 516232 441594 516364 441600
rect 516140 441584 516192 441590
rect 516244 441586 516364 441594
rect 516140 441526 516192 441532
rect 516152 440609 516180 441526
rect 516138 440600 516194 440609
rect 516138 440535 516194 440544
rect 513746 440328 513802 440337
rect 513746 440263 513748 440272
rect 513800 440263 513802 440272
rect 513748 440234 513800 440240
rect 516138 438968 516194 438977
rect 516138 438903 516140 438912
rect 516192 438903 516194 438912
rect 516140 438874 516192 438880
rect 516230 438424 516286 438433
rect 516230 438359 516286 438368
rect 516138 437880 516194 437889
rect 516138 437815 516194 437824
rect 516152 437510 516180 437815
rect 516244 437578 516272 438359
rect 516232 437572 516284 437578
rect 516232 437514 516284 437520
rect 516140 437504 516192 437510
rect 516140 437446 516192 437452
rect 516230 437336 516286 437345
rect 516230 437271 516286 437280
rect 516244 436286 516272 437271
rect 516232 436280 516284 436286
rect 516138 436248 516194 436257
rect 516232 436222 516284 436228
rect 516138 436183 516194 436192
rect 516152 436150 516180 436183
rect 516140 436144 516192 436150
rect 516140 436086 516192 436092
rect 516230 435704 516286 435713
rect 516230 435639 516286 435648
rect 516138 435160 516194 435169
rect 516138 435095 516194 435104
rect 516152 434858 516180 435095
rect 516140 434852 516192 434858
rect 516140 434794 516192 434800
rect 516244 434790 516272 435639
rect 516232 434784 516284 434790
rect 516232 434726 516284 434732
rect 516230 434072 516286 434081
rect 516230 434007 516286 434016
rect 516138 433528 516194 433537
rect 516138 433463 516140 433472
rect 516192 433463 516194 433472
rect 516140 433434 516192 433440
rect 516244 433362 516272 434007
rect 516232 433356 516284 433362
rect 516232 433298 516284 433304
rect 513470 432304 513526 432313
rect 513470 432239 513526 432248
rect 516336 432154 516364 441586
rect 516060 432126 516364 432154
rect 516060 431954 516088 432126
rect 516230 432032 516286 432041
rect 516230 431967 516286 431976
rect 516060 431926 516180 431954
rect 513378 430672 513434 430681
rect 513378 430607 513434 430616
rect 516152 426601 516180 431926
rect 516244 431497 516272 431967
rect 516230 431488 516286 431497
rect 516230 431423 516286 431432
rect 516428 430953 516456 460158
rect 516600 442264 516652 442270
rect 516600 442206 516652 442212
rect 516508 441720 516560 441726
rect 516508 441662 516560 441668
rect 516520 436898 516548 441662
rect 516508 436892 516560 436898
rect 516508 436834 516560 436840
rect 516506 436792 516562 436801
rect 516506 436727 516562 436736
rect 516520 436218 516548 436727
rect 516508 436212 516560 436218
rect 516508 436154 516560 436160
rect 516506 434616 516562 434625
rect 516506 434551 516562 434560
rect 516520 433430 516548 434551
rect 516508 433424 516560 433430
rect 516508 433366 516560 433372
rect 516506 432984 516562 432993
rect 516506 432919 516562 432928
rect 516520 432070 516548 432919
rect 516508 432064 516560 432070
rect 516508 432006 516560 432012
rect 516612 431954 516640 442206
rect 516692 441924 516744 441930
rect 516692 441866 516744 441872
rect 516520 431926 516640 431954
rect 516414 430944 516470 430953
rect 516414 430879 516470 430888
rect 516414 429856 516470 429865
rect 516414 429791 516470 429800
rect 516428 429162 516456 429791
rect 516520 429321 516548 431926
rect 516506 429312 516562 429321
rect 516506 429247 516562 429256
rect 516428 429134 516548 429162
rect 516414 428768 516470 428777
rect 516414 428703 516470 428712
rect 516138 426592 516194 426601
rect 516138 426527 516194 426536
rect 516322 426048 516378 426057
rect 516322 425983 516378 425992
rect 516138 424960 516194 424969
rect 516138 424895 516194 424904
rect 516152 424590 516180 424895
rect 516140 424584 516192 424590
rect 516140 424526 516192 424532
rect 516140 424448 516192 424454
rect 516138 424416 516140 424425
rect 516192 424416 516194 424425
rect 516138 424351 516194 424360
rect 516232 424380 516284 424386
rect 516232 424322 516284 424328
rect 516244 423881 516272 424322
rect 516230 423872 516286 423881
rect 516230 423807 516286 423816
rect 516336 423722 516364 425983
rect 516244 423694 516364 423722
rect 516138 423328 516194 423337
rect 516138 423263 516194 423272
rect 516152 422550 516180 423263
rect 516140 422544 516192 422550
rect 516140 422486 516192 422492
rect 516140 422408 516192 422414
rect 516140 422350 516192 422356
rect 504560 412134 504942 412162
rect 500224 412072 500276 412078
rect 500224 412014 500276 412020
rect 497464 412004 497516 412010
rect 497464 411946 497516 411952
rect 497476 358766 497504 411946
rect 497464 358760 497516 358766
rect 497464 358702 497516 358708
rect 500236 357406 500264 412014
rect 504560 409766 504588 412134
rect 516152 412078 516180 422350
rect 516244 412622 516272 423694
rect 516322 422784 516378 422793
rect 516322 422719 516378 422728
rect 516336 422346 516364 422719
rect 516428 422482 516456 428703
rect 516416 422476 516468 422482
rect 516416 422418 516468 422424
rect 516520 422362 516548 429134
rect 516704 427145 516732 441866
rect 516888 439142 516916 494935
rect 517256 493921 517284 560351
rect 517440 495009 517468 560895
rect 517532 554810 517560 574926
rect 520372 568948 520424 568954
rect 520372 568890 520424 568896
rect 517702 568440 517758 568449
rect 517702 568375 517758 568384
rect 517610 565856 517666 565865
rect 517610 565791 517666 565800
rect 517520 554804 517572 554810
rect 517520 554746 517572 554752
rect 517624 505442 517652 565791
rect 517716 511193 517744 568375
rect 519360 567316 519412 567322
rect 519360 567258 519412 567264
rect 519268 564528 519320 564534
rect 519268 564470 519320 564476
rect 518992 563304 519044 563310
rect 518992 563246 519044 563252
rect 517796 563100 517848 563106
rect 517796 563042 517848 563048
rect 517808 520946 517836 563042
rect 517888 562012 517940 562018
rect 517888 561954 517940 561960
rect 517900 526454 517928 561954
rect 517980 561468 518032 561474
rect 517980 561410 518032 561416
rect 517888 526448 517940 526454
rect 517888 526390 517940 526396
rect 517796 520940 517848 520946
rect 517796 520882 517848 520888
rect 517702 511184 517758 511193
rect 517702 511119 517758 511128
rect 517716 510678 517744 511119
rect 517704 510672 517756 510678
rect 517704 510614 517756 510620
rect 517612 505436 517664 505442
rect 517612 505378 517664 505384
rect 517808 500546 517836 520882
rect 517796 500540 517848 500546
rect 517796 500482 517848 500488
rect 517900 498166 517928 526390
rect 517888 498160 517940 498166
rect 517888 498102 517940 498108
rect 517992 495514 518020 561410
rect 518164 514072 518216 514078
rect 518164 514014 518216 514020
rect 517520 495508 517572 495514
rect 517520 495450 517572 495456
rect 517980 495508 518032 495514
rect 517980 495450 518032 495456
rect 517426 495000 517482 495009
rect 517426 494935 517482 494944
rect 517242 493912 517298 493921
rect 517242 493847 517298 493856
rect 517244 488504 517296 488510
rect 517244 488446 517296 488452
rect 517256 488073 517284 488446
rect 517242 488064 517298 488073
rect 517242 487999 517298 488008
rect 516968 441856 517020 441862
rect 516968 441798 517020 441804
rect 516876 439136 516928 439142
rect 516876 439078 516928 439084
rect 516876 436892 516928 436898
rect 516876 436834 516928 436840
rect 516782 432440 516838 432449
rect 516782 432375 516838 432384
rect 516796 432002 516824 432375
rect 516888 432041 516916 436834
rect 516874 432032 516930 432041
rect 516784 431996 516836 432002
rect 516874 431967 516930 431976
rect 516784 431938 516836 431944
rect 516782 428224 516838 428233
rect 516782 428159 516838 428168
rect 516690 427136 516746 427145
rect 516690 427071 516746 427080
rect 516796 426986 516824 428159
rect 516980 427689 517008 441798
rect 517058 441688 517114 441697
rect 517058 441623 517114 441632
rect 516966 427680 517022 427689
rect 516966 427615 517022 427624
rect 516324 422340 516376 422346
rect 516324 422282 516376 422288
rect 516428 422334 516548 422362
rect 516704 426958 516824 426986
rect 516322 422240 516378 422249
rect 516322 422175 516378 422184
rect 516336 421938 516364 422175
rect 516324 421932 516376 421938
rect 516324 421874 516376 421880
rect 516322 421832 516378 421841
rect 516322 421767 516378 421776
rect 516336 421598 516364 421767
rect 516324 421592 516376 421598
rect 516324 421534 516376 421540
rect 516322 421288 516378 421297
rect 516322 421223 516378 421232
rect 516336 421190 516364 421223
rect 516324 421184 516376 421190
rect 516324 421126 516376 421132
rect 516322 420744 516378 420753
rect 516322 420679 516378 420688
rect 516336 419830 516364 420679
rect 516324 419824 516376 419830
rect 516324 419766 516376 419772
rect 516322 418568 516378 418577
rect 516322 418503 516324 418512
rect 516376 418503 516378 418512
rect 516324 418474 516376 418480
rect 516322 418024 516378 418033
rect 516322 417959 516378 417968
rect 516336 417450 516364 417959
rect 516324 417444 516376 417450
rect 516324 417386 516376 417392
rect 516322 415848 516378 415857
rect 516322 415783 516324 415792
rect 516376 415783 516378 415792
rect 516324 415754 516376 415760
rect 516322 414760 516378 414769
rect 516322 414695 516324 414704
rect 516376 414695 516378 414704
rect 516324 414666 516376 414672
rect 516322 414216 516378 414225
rect 516322 414151 516378 414160
rect 516336 414118 516364 414151
rect 516324 414112 516376 414118
rect 516324 414054 516376 414060
rect 516324 413296 516376 413302
rect 516324 413238 516376 413244
rect 516336 413137 516364 413238
rect 516322 413128 516378 413137
rect 516322 413063 516378 413072
rect 516232 412616 516284 412622
rect 516232 412558 516284 412564
rect 516322 412584 516378 412593
rect 516322 412519 516324 412528
rect 516376 412519 516378 412528
rect 516324 412490 516376 412496
rect 516140 412072 516192 412078
rect 506874 411998 506980 412026
rect 508898 411998 509004 412026
rect 510922 411998 511028 412026
rect 512946 411998 513052 412026
rect 516140 412014 516192 412020
rect 516428 412010 516456 422334
rect 516506 419112 516562 419121
rect 516506 419047 516562 419056
rect 516520 418606 516548 419047
rect 516508 418600 516560 418606
rect 516508 418542 516560 418548
rect 516600 417376 516652 417382
rect 516600 417318 516652 417324
rect 516612 416945 516640 417318
rect 516598 416936 516654 416945
rect 516598 416871 516654 416880
rect 516506 416392 516562 416401
rect 516506 416327 516562 416336
rect 516520 415478 516548 416327
rect 516508 415472 516560 415478
rect 516508 415414 516560 415420
rect 516506 415304 516562 415313
rect 516506 415239 516562 415248
rect 516520 414050 516548 415239
rect 516508 414044 516560 414050
rect 516508 413986 516560 413992
rect 516704 412634 516732 426958
rect 516784 425740 516836 425746
rect 516784 425682 516836 425688
rect 516796 425513 516824 425682
rect 516782 425504 516838 425513
rect 516782 425439 516838 425448
rect 516784 420232 516836 420238
rect 516782 420200 516784 420209
rect 516836 420200 516838 420209
rect 516782 420135 516838 420144
rect 516784 420028 516836 420034
rect 516784 419970 516836 419976
rect 516796 419665 516824 419970
rect 516782 419656 516838 419665
rect 516782 419591 516838 419600
rect 516782 413672 516838 413681
rect 516782 413607 516838 413616
rect 516796 412690 516824 413607
rect 516520 412606 516732 412634
rect 516784 412684 516836 412690
rect 516784 412626 516836 412632
rect 504548 409760 504600 409766
rect 504548 409702 504600 409708
rect 501604 409148 501656 409154
rect 501604 409090 501656 409096
rect 500224 357400 500276 357406
rect 500224 357342 500276 357348
rect 494060 304768 494112 304774
rect 494060 304710 494112 304716
rect 471060 269068 471112 269074
rect 471060 269010 471112 269016
rect 471244 269068 471296 269074
rect 471244 269010 471296 269016
rect 471072 268530 471100 269010
rect 486424 268592 486476 268598
rect 486424 268534 486476 268540
rect 471060 268524 471112 268530
rect 471060 268466 471112 268472
rect 476764 268524 476816 268530
rect 476764 268466 476816 268472
rect 457444 268456 457496 268462
rect 457444 268398 457496 268404
rect 456064 225004 456116 225010
rect 456064 224946 456116 224952
rect 456076 222154 456104 224946
rect 454684 222148 454736 222154
rect 454684 222090 454736 222096
rect 456064 222148 456116 222154
rect 456064 222090 456116 222096
rect 450544 209160 450596 209166
rect 450544 209102 450596 209108
rect 449256 208344 449308 208350
rect 449256 208286 449308 208292
rect 448152 205896 448204 205902
rect 448152 205838 448204 205844
rect 447968 205624 448020 205630
rect 447968 205566 448020 205572
rect 447232 202836 447284 202842
rect 447232 202778 447284 202784
rect 447876 202836 447928 202842
rect 447876 202778 447928 202784
rect 447244 201550 447272 202778
rect 447232 201544 447284 201550
rect 447232 201486 447284 201492
rect 447140 197260 447192 197266
rect 447140 197202 447192 197208
rect 447152 196722 447180 197202
rect 447140 196716 447192 196722
rect 447140 196658 447192 196664
rect 446496 196104 446548 196110
rect 446496 196046 446548 196052
rect 446048 190426 446444 190454
rect 446416 189106 446444 190426
rect 446404 189100 446456 189106
rect 446404 189042 446456 189048
rect 445772 180766 445892 180794
rect 445300 163804 445352 163810
rect 445300 163746 445352 163752
rect 445208 162852 445260 162858
rect 445208 162794 445260 162800
rect 445208 156664 445260 156670
rect 445208 156606 445260 156612
rect 445220 154562 445248 156606
rect 445208 154556 445260 154562
rect 445208 154498 445260 154504
rect 445116 153740 445168 153746
rect 445116 153682 445168 153688
rect 445128 143177 445156 153682
rect 445114 143168 445170 143177
rect 445114 143103 445170 143112
rect 445220 141953 445248 154498
rect 445312 153814 445340 163746
rect 445576 154488 445628 154494
rect 445576 154430 445628 154436
rect 445300 153808 445352 153814
rect 445300 153750 445352 153756
rect 445312 148889 445340 153750
rect 445588 153474 445616 154430
rect 445576 153468 445628 153474
rect 445576 153410 445628 153416
rect 445298 148880 445354 148889
rect 445298 148815 445354 148824
rect 445206 141944 445262 141953
rect 445206 141879 445262 141888
rect 445588 139641 445616 153410
rect 445668 152516 445720 152522
rect 445668 152458 445720 152464
rect 445680 152425 445708 152458
rect 445666 152416 445722 152425
rect 445666 152351 445722 152360
rect 445574 139632 445630 139641
rect 445574 139567 445630 139576
rect 445298 137320 445354 137329
rect 445298 137255 445354 137264
rect 445312 136678 445340 137255
rect 445300 136672 445352 136678
rect 445300 136614 445352 136620
rect 445024 135312 445076 135318
rect 445024 135254 445076 135260
rect 445668 135312 445720 135318
rect 445668 135254 445720 135260
rect 445116 133952 445168 133958
rect 445680 133929 445708 135254
rect 445116 133894 445168 133900
rect 445666 133920 445722 133929
rect 445128 132705 445156 133894
rect 445666 133855 445722 133864
rect 445114 132696 445170 132705
rect 445114 132631 445170 132640
rect 445116 132524 445168 132530
rect 445116 132466 445168 132472
rect 445128 132161 445156 132466
rect 445114 132152 445170 132161
rect 445114 132087 445170 132096
rect 443368 127628 443420 127634
rect 443368 127570 443420 127576
rect 444932 127628 444984 127634
rect 444932 127570 444984 127576
rect 443380 125934 443408 127570
rect 444932 126336 444984 126342
rect 444932 126278 444984 126284
rect 444840 126268 444892 126274
rect 444840 126210 444892 126216
rect 443368 125928 443420 125934
rect 443368 125870 443420 125876
rect 443092 125452 443144 125458
rect 443092 125394 443144 125400
rect 444852 125390 444880 126210
rect 444944 125526 444972 126278
rect 444932 125520 444984 125526
rect 444932 125462 444984 125468
rect 442080 125384 442132 125390
rect 442080 125326 442132 125332
rect 444840 125384 444892 125390
rect 444840 125326 444892 125332
rect 445772 125254 445800 180766
rect 445852 160880 445904 160886
rect 445852 160822 445904 160828
rect 445864 160750 445892 160822
rect 445852 160744 445904 160750
rect 445852 160686 445904 160692
rect 445864 138553 445892 160686
rect 445942 156496 445998 156505
rect 445942 156431 445998 156440
rect 445956 156097 445984 156431
rect 445942 156088 445998 156097
rect 445942 156023 445998 156032
rect 445956 151201 445984 156023
rect 446416 153950 446444 189042
rect 446508 160886 446536 196046
rect 446496 160880 446548 160886
rect 446496 160822 446548 160828
rect 446404 153944 446456 153950
rect 446404 153886 446456 153892
rect 445942 151192 445998 151201
rect 445942 151127 445998 151136
rect 445850 138544 445906 138553
rect 445850 138479 445906 138488
rect 445864 138038 445892 138479
rect 445852 138032 445904 138038
rect 445852 137974 445904 137980
rect 446404 138032 446456 138038
rect 446404 137974 446456 137980
rect 445760 125248 445812 125254
rect 445760 125190 445812 125196
rect 446416 124982 446444 137974
rect 447244 135930 447272 201486
rect 450556 152522 450584 209102
rect 454696 207670 454724 222090
rect 457456 212362 457484 268398
rect 464344 225072 464396 225078
rect 464344 225014 464396 225020
rect 461584 223916 461636 223922
rect 461584 223858 461636 223864
rect 457444 212356 457496 212362
rect 457444 212298 457496 212304
rect 461596 209166 461624 223858
rect 461584 209160 461636 209166
rect 461584 209102 461636 209108
rect 464356 209098 464384 225014
rect 475384 218136 475436 218142
rect 475384 218078 475436 218084
rect 471244 217320 471296 217326
rect 471244 217262 471296 217268
rect 468484 215960 468536 215966
rect 468484 215902 468536 215908
rect 464344 209092 464396 209098
rect 464344 209034 464396 209040
rect 454684 207664 454736 207670
rect 454684 207606 454736 207612
rect 466920 196852 466972 196858
rect 466920 196794 466972 196800
rect 457444 196716 457496 196722
rect 457444 196658 457496 196664
rect 450544 152516 450596 152522
rect 450544 152458 450596 152464
rect 447232 135924 447284 135930
rect 447232 135866 447284 135872
rect 457456 126274 457484 196658
rect 460204 196648 460256 196654
rect 460204 196590 460256 196596
rect 460216 154562 460244 196590
rect 466932 196042 466960 196794
rect 466920 196036 466972 196042
rect 466920 195978 466972 195984
rect 466932 190454 466960 195978
rect 466932 190426 467144 190454
rect 459744 154556 459796 154562
rect 459744 154498 459796 154504
rect 460204 154556 460256 154562
rect 460204 154498 460256 154504
rect 459756 154018 459784 154498
rect 459744 154012 459796 154018
rect 459744 153954 459796 153960
rect 467116 126342 467144 190426
rect 468496 155242 468524 215902
rect 468484 155236 468536 155242
rect 468484 155178 468536 155184
rect 471256 152590 471284 217262
rect 472624 216708 472676 216714
rect 472624 216650 472676 216656
rect 472636 152658 472664 216650
rect 475396 152726 475424 218078
rect 476776 212430 476804 268466
rect 483664 222352 483716 222358
rect 483664 222294 483716 222300
rect 482284 220924 482336 220930
rect 482284 220866 482336 220872
rect 479524 219632 479576 219638
rect 479524 219574 479576 219580
rect 476764 212424 476816 212430
rect 476764 212366 476816 212372
rect 476488 198008 476540 198014
rect 476488 197950 476540 197956
rect 476500 197402 476528 197950
rect 476488 197396 476540 197402
rect 476488 197338 476540 197344
rect 476764 197396 476816 197402
rect 476764 197338 476816 197344
rect 475384 152720 475436 152726
rect 475384 152662 475436 152668
rect 472624 152652 472676 152658
rect 472624 152594 472676 152600
rect 471244 152584 471296 152590
rect 471244 152526 471296 152532
rect 476776 129062 476804 197338
rect 479536 153202 479564 219574
rect 482296 154086 482324 220866
rect 482284 154080 482336 154086
rect 482284 154022 482336 154028
rect 483676 153921 483704 222294
rect 485044 222216 485096 222222
rect 485044 222158 485096 222164
rect 485056 154154 485084 222158
rect 486436 212498 486464 268534
rect 489184 222284 489236 222290
rect 489184 222226 489236 222232
rect 486424 212492 486476 212498
rect 486424 212434 486476 212440
rect 489196 154222 489224 222226
rect 490564 220856 490616 220862
rect 490564 220798 490616 220804
rect 489184 154216 489236 154222
rect 489184 154158 489236 154164
rect 485044 154148 485096 154154
rect 485044 154090 485096 154096
rect 483662 153912 483718 153921
rect 483662 153847 483718 153856
rect 479524 153196 479576 153202
rect 479524 153138 479576 153144
rect 490576 152794 490604 220798
rect 493324 219564 493376 219570
rect 493324 219506 493376 219512
rect 493336 153134 493364 219506
rect 494704 219496 494756 219502
rect 494704 219438 494756 219444
rect 493324 153128 493376 153134
rect 493324 153070 493376 153076
rect 494716 152862 494744 219438
rect 497464 218068 497516 218074
rect 497464 218010 497516 218016
rect 497476 152930 497504 218010
rect 497464 152924 497516 152930
rect 497464 152866 497516 152872
rect 494704 152856 494756 152862
rect 494704 152798 494756 152804
rect 490564 152788 490616 152794
rect 490564 152730 490616 152736
rect 497464 136672 497516 136678
rect 497464 136614 497516 136620
rect 490564 134020 490616 134026
rect 490564 133962 490616 133968
rect 476764 129056 476816 129062
rect 476764 128998 476816 129004
rect 467104 126336 467156 126342
rect 467104 126278 467156 126284
rect 457444 126268 457496 126274
rect 457444 126210 457496 126216
rect 446404 124976 446456 124982
rect 446404 124918 446456 124924
rect 490576 124914 490604 133962
rect 493968 126336 494020 126342
rect 493968 126278 494020 126284
rect 493980 125186 494008 126278
rect 494704 126268 494756 126274
rect 494704 126210 494756 126216
rect 493968 125180 494020 125186
rect 493968 125122 494020 125128
rect 494716 125118 494744 126210
rect 494704 125112 494756 125118
rect 494704 125054 494756 125060
rect 490564 124908 490616 124914
rect 490564 124850 490616 124856
rect 497476 124846 497504 136614
rect 500224 135924 500276 135930
rect 500224 135866 500276 135872
rect 500236 125050 500264 135866
rect 500224 125044 500276 125050
rect 500224 124986 500276 124992
rect 497464 124840 497516 124846
rect 497464 124782 497516 124788
rect 441712 122664 441764 122670
rect 441712 122606 441764 122612
rect 438860 122596 438912 122602
rect 438860 122538 438912 122544
rect 431224 99544 431276 99550
rect 431224 99486 431276 99492
rect 501616 99482 501644 409090
rect 506952 393314 506980 411998
rect 508976 409834 509004 411998
rect 508964 409828 509016 409834
rect 508964 409770 509016 409776
rect 511000 409154 511028 411998
rect 513024 409698 513052 411998
rect 516416 412004 516468 412010
rect 516416 411946 516468 411952
rect 516520 411942 516548 412606
rect 516508 411936 516560 411942
rect 516508 411878 516560 411884
rect 513378 411632 513434 411641
rect 513378 411567 513434 411576
rect 513392 411330 513420 411567
rect 513380 411324 513432 411330
rect 513380 411266 513432 411272
rect 513012 409692 513064 409698
rect 513012 409634 513064 409640
rect 510988 409148 511040 409154
rect 510988 409090 511040 409096
rect 506492 393286 506980 393314
rect 506492 370530 506520 393286
rect 516600 377460 516652 377466
rect 516600 377402 516652 377408
rect 516612 376786 516640 377402
rect 516416 376780 516468 376786
rect 516416 376722 516468 376728
rect 516600 376780 516652 376786
rect 516600 376722 516652 376728
rect 516140 371748 516192 371754
rect 516140 371690 516192 371696
rect 516152 371278 516180 371690
rect 516140 371272 516192 371278
rect 516140 371214 516192 371220
rect 506480 370524 506532 370530
rect 506480 370466 506532 370472
rect 513380 370524 513432 370530
rect 513380 370466 513432 370472
rect 502984 367872 503036 367878
rect 502984 367814 503036 367820
rect 502996 352578 503024 367814
rect 502984 352572 503036 352578
rect 502984 352514 503036 352520
rect 513392 345014 513420 370466
rect 516152 370002 516180 371214
rect 516152 369974 516272 370002
rect 516140 369844 516192 369850
rect 516140 369786 516192 369792
rect 516152 369481 516180 369786
rect 516138 369472 516194 369481
rect 516138 369407 516194 369416
rect 513746 369200 513802 369209
rect 513746 369135 513748 369144
rect 513800 369135 513802 369144
rect 513748 369106 513800 369112
rect 516140 368416 516192 368422
rect 516138 368384 516140 368393
rect 516192 368384 516194 368393
rect 516138 368319 516194 368328
rect 513654 367976 513710 367985
rect 513654 367911 513656 367920
rect 513708 367911 513710 367920
rect 513656 367882 513708 367888
rect 513748 367872 513800 367878
rect 513748 367814 513800 367820
rect 513760 367713 513788 367814
rect 516140 367804 516192 367810
rect 516140 367746 516192 367752
rect 513746 367704 513802 367713
rect 513746 367639 513802 367648
rect 516152 367169 516180 367746
rect 516138 367160 516194 367169
rect 516138 367095 516194 367104
rect 516244 364857 516272 369974
rect 516428 366081 516456 376722
rect 516414 366072 516470 366081
rect 516414 366007 516470 366016
rect 516230 364848 516286 364857
rect 516230 364783 516286 364792
rect 516138 363760 516194 363769
rect 516138 363695 516194 363704
rect 516152 363662 516180 363695
rect 516140 363656 516192 363662
rect 516140 363598 516192 363604
rect 516140 362704 516192 362710
rect 516140 362646 516192 362652
rect 516152 362545 516180 362646
rect 516138 362536 516194 362545
rect 516138 362471 516194 362480
rect 516782 361448 516838 361457
rect 516782 361383 516838 361392
rect 516796 360874 516824 361383
rect 516784 360868 516836 360874
rect 516784 360810 516836 360816
rect 516140 360732 516192 360738
rect 516140 360674 516192 360680
rect 516152 360233 516180 360674
rect 516138 360224 516194 360233
rect 516138 360159 516194 360168
rect 516140 359168 516192 359174
rect 516138 359136 516140 359145
rect 516192 359136 516194 359145
rect 516138 359071 516194 359080
rect 516140 357944 516192 357950
rect 516138 357912 516140 357921
rect 516192 357912 516194 357921
rect 516138 357847 516194 357856
rect 516416 357400 516468 357406
rect 516416 357342 516468 357348
rect 516428 356833 516456 357342
rect 516414 356824 516470 356833
rect 516414 356759 516470 356768
rect 516140 355632 516192 355638
rect 516138 355600 516140 355609
rect 516192 355600 516194 355609
rect 516138 355535 516194 355544
rect 516140 354544 516192 354550
rect 516138 354512 516140 354521
rect 516192 354512 516194 354521
rect 516138 354447 516194 354456
rect 516140 351892 516192 351898
rect 516140 351834 516192 351840
rect 516152 350985 516180 351834
rect 516138 350976 516194 350985
rect 516138 350911 516194 350920
rect 516140 348832 516192 348838
rect 516140 348774 516192 348780
rect 516152 348673 516180 348774
rect 516138 348664 516194 348673
rect 516138 348599 516194 348608
rect 516138 347576 516194 347585
rect 516138 347511 516194 347520
rect 516152 347070 516180 347511
rect 516140 347064 516192 347070
rect 516140 347006 516192 347012
rect 516232 346384 516284 346390
rect 516138 346352 516194 346361
rect 516232 346326 516284 346332
rect 516138 346287 516140 346296
rect 516192 346287 516194 346296
rect 516140 346258 516192 346264
rect 516244 345273 516272 346326
rect 516230 345264 516286 345273
rect 516230 345199 516286 345208
rect 513392 344986 513512 345014
rect 513378 340912 513434 340921
rect 513378 340847 513434 340856
rect 513392 340814 513420 340847
rect 513380 340808 513432 340814
rect 513380 340750 513432 340756
rect 503732 340054 504942 340082
rect 503732 266354 503760 340054
rect 506860 338094 506888 340068
rect 507872 340054 508898 340082
rect 506848 338088 506900 338094
rect 506848 338030 506900 338036
rect 507768 338088 507820 338094
rect 507768 338030 507820 338036
rect 507780 298518 507808 338030
rect 507768 298512 507820 298518
rect 507768 298454 507820 298460
rect 507872 297906 507900 340054
rect 510908 337414 510936 340068
rect 512932 337754 512960 340068
rect 513484 338094 513512 344986
rect 516140 344344 516192 344350
rect 516140 344286 516192 344292
rect 516152 344049 516180 344286
rect 516138 344040 516194 344049
rect 516138 343975 516194 343984
rect 514760 343596 514812 343602
rect 514760 343538 514812 343544
rect 514772 342961 514800 343538
rect 514758 342952 514814 342961
rect 514758 342887 514814 342896
rect 514772 342106 514800 342887
rect 514760 342100 514812 342106
rect 514760 342042 514812 342048
rect 516140 341760 516192 341766
rect 516138 341728 516140 341737
rect 516192 341728 516194 341737
rect 516138 341663 516194 341672
rect 516428 340882 516456 356759
rect 516598 349888 516654 349897
rect 516598 349823 516600 349832
rect 516652 349823 516654 349832
rect 516600 349794 516652 349800
rect 516416 340876 516468 340882
rect 516416 340818 516468 340824
rect 513472 338088 513524 338094
rect 513472 338030 513524 338036
rect 512920 337748 512972 337754
rect 512920 337690 512972 337696
rect 514760 337748 514812 337754
rect 514760 337690 514812 337696
rect 510896 337408 510948 337414
rect 510896 337350 510948 337356
rect 514208 298512 514260 298518
rect 514208 298454 514260 298460
rect 507860 297900 507912 297906
rect 507860 297842 507912 297848
rect 513748 297900 513800 297906
rect 513748 297842 513800 297848
rect 513378 297528 513434 297537
rect 513378 297463 513434 297472
rect 513392 297430 513420 297463
rect 513380 297424 513432 297430
rect 513380 297366 513432 297372
rect 513288 297220 513340 297226
rect 513288 297162 513340 297168
rect 513300 296290 513328 297162
rect 513378 296848 513434 296857
rect 513378 296783 513434 296792
rect 513392 296750 513420 296783
rect 513380 296744 513432 296750
rect 513380 296686 513432 296692
rect 513380 296608 513432 296614
rect 513380 296550 513432 296556
rect 513392 296449 513420 296550
rect 513472 296472 513524 296478
rect 513378 296440 513434 296449
rect 513472 296414 513524 296420
rect 513378 296375 513434 296384
rect 513300 296262 513420 296290
rect 513392 286249 513420 296262
rect 513484 295905 513512 296414
rect 513562 296304 513618 296313
rect 513562 296239 513618 296248
rect 513470 295896 513526 295905
rect 513576 295866 513604 296239
rect 513470 295831 513526 295840
rect 513564 295860 513616 295866
rect 513564 295802 513616 295808
rect 513760 295746 513788 297842
rect 514116 297288 514168 297294
rect 514116 297230 514168 297236
rect 513932 297152 513984 297158
rect 513932 297094 513984 297100
rect 513840 297084 513892 297090
rect 513840 297026 513892 297032
rect 513484 295718 513788 295746
rect 513378 286240 513434 286249
rect 513378 286175 513434 286184
rect 513380 269068 513432 269074
rect 513380 269010 513432 269016
rect 513288 269000 513340 269006
rect 513288 268942 513340 268948
rect 513300 268682 513328 268942
rect 512946 268668 513328 268682
rect 512932 268654 513328 268668
rect 504928 266354 504956 268124
rect 506860 266354 506888 268124
rect 503720 266348 503772 266354
rect 503720 266290 503772 266296
rect 504916 266348 504968 266354
rect 504916 266290 504968 266296
rect 506848 266348 506900 266354
rect 506848 266290 506900 266296
rect 507768 266348 507820 266354
rect 507768 266290 507820 266296
rect 503732 265742 503760 266290
rect 503720 265736 503772 265742
rect 503720 265678 503772 265684
rect 502984 264988 503036 264994
rect 502984 264930 503036 264936
rect 501604 99476 501656 99482
rect 501604 99418 501656 99424
rect 502996 99414 503024 264930
rect 503732 209774 503760 265678
rect 507780 225622 507808 266290
rect 508884 266286 508912 268124
rect 508872 266280 508924 266286
rect 508872 266222 508924 266228
rect 509148 266280 509200 266286
rect 509148 266222 509200 266228
rect 509160 225690 509188 266222
rect 510908 264994 510936 268124
rect 512932 267734 512960 268654
rect 513392 268433 513420 269010
rect 513378 268424 513434 268433
rect 513378 268359 513434 268368
rect 512656 267706 512960 267734
rect 512656 265674 512684 267706
rect 513484 266286 513512 295718
rect 513852 295610 513880 297026
rect 513576 295582 513880 295610
rect 513576 286793 513604 295582
rect 513656 295520 513708 295526
rect 513944 295474 513972 297094
rect 513656 295462 513708 295468
rect 513668 287881 513696 295462
rect 513852 295446 513972 295474
rect 513748 291916 513800 291922
rect 513748 291858 513800 291864
rect 513654 287872 513710 287881
rect 513654 287807 513710 287816
rect 513562 286784 513618 286793
rect 513562 286719 513618 286728
rect 513760 266354 513788 291858
rect 513852 286793 513880 295446
rect 514128 295202 514156 297230
rect 513944 295174 514156 295202
rect 513944 288289 513972 295174
rect 514220 292574 514248 298454
rect 514036 292546 514248 292574
rect 514036 291922 514064 292546
rect 514024 291916 514076 291922
rect 514024 291858 514076 291864
rect 513930 288280 513986 288289
rect 513930 288215 513986 288224
rect 513838 286784 513894 286793
rect 513838 286719 513894 286728
rect 514772 269006 514800 337690
rect 517072 306374 517100 441623
rect 517334 441144 517390 441153
rect 517334 441079 517390 441088
rect 517242 440056 517298 440065
rect 517242 439991 517298 440000
rect 516980 306346 517100 306374
rect 515404 299736 515456 299742
rect 515404 299678 515456 299684
rect 514760 269000 514812 269006
rect 514760 268942 514812 268948
rect 513748 266348 513800 266354
rect 513748 266290 513800 266296
rect 513472 266280 513524 266286
rect 513472 266222 513524 266228
rect 512644 265668 512696 265674
rect 512644 265610 512696 265616
rect 510896 264988 510948 264994
rect 510896 264930 510948 264936
rect 509148 225684 509200 225690
rect 509148 225626 509200 225632
rect 512656 225622 512684 265610
rect 514852 225684 514904 225690
rect 514852 225626 514904 225632
rect 507768 225616 507820 225622
rect 507768 225558 507820 225564
rect 512644 225616 512696 225622
rect 512644 225558 512696 225564
rect 514760 225548 514812 225554
rect 514760 225490 514812 225496
rect 513748 225072 513800 225078
rect 513746 225040 513748 225049
rect 513800 225040 513802 225049
rect 513380 225004 513432 225010
rect 513746 224975 513802 224984
rect 513380 224946 513432 224952
rect 513392 221921 513420 224946
rect 513746 223952 513802 223961
rect 513746 223887 513748 223896
rect 513800 223887 513802 223896
rect 513748 223858 513800 223864
rect 513378 221912 513434 221921
rect 513378 221847 513434 221856
rect 503732 209746 504496 209774
rect 504468 196738 504496 209746
rect 514668 201272 514720 201278
rect 514666 201240 514668 201249
rect 514720 201240 514722 201249
rect 514666 201175 514722 201184
rect 513562 200832 513618 200841
rect 513562 200767 513618 200776
rect 513378 199472 513434 199481
rect 513378 199407 513434 199416
rect 513392 198014 513420 199407
rect 513576 198082 513604 200767
rect 514208 200116 514260 200122
rect 514208 200058 514260 200064
rect 514116 200048 514168 200054
rect 514114 200016 514116 200025
rect 514168 200016 514170 200025
rect 514114 199951 514170 199960
rect 514220 198937 514248 200058
rect 514206 198928 514262 198937
rect 514206 198863 514262 198872
rect 514116 198688 514168 198694
rect 514116 198630 514168 198636
rect 513564 198076 513616 198082
rect 513564 198018 513616 198024
rect 513380 198008 513432 198014
rect 513380 197950 513432 197956
rect 514128 197713 514156 198630
rect 514114 197704 514170 197713
rect 514114 197639 514170 197648
rect 513288 197328 513340 197334
rect 513288 197270 513340 197276
rect 513300 196738 513328 197270
rect 504468 196710 504942 196738
rect 512946 196710 513328 196738
rect 514128 196722 514156 197639
rect 514220 196858 514248 198863
rect 514208 196852 514260 196858
rect 514208 196794 514260 196800
rect 514116 196716 514168 196722
rect 514116 196658 514168 196664
rect 506860 194478 506888 196044
rect 506848 194472 506900 194478
rect 506848 194414 506900 194420
rect 507768 194472 507820 194478
rect 507768 194414 507820 194420
rect 507780 155310 507808 194414
rect 508884 194410 508912 196044
rect 510908 194546 510936 196044
rect 510896 194540 510948 194546
rect 510896 194482 510948 194488
rect 514772 194478 514800 225490
rect 514760 194472 514812 194478
rect 514760 194414 514812 194420
rect 514864 194410 514892 225626
rect 514944 225616 514996 225622
rect 514944 225558 514996 225564
rect 514956 197334 514984 225558
rect 515416 206854 515444 299678
rect 516784 298852 516836 298858
rect 516784 298794 516836 298800
rect 516600 298784 516652 298790
rect 516600 298726 516652 298732
rect 516508 298376 516560 298382
rect 516508 298318 516560 298324
rect 516324 297560 516376 297566
rect 516324 297502 516376 297508
rect 516232 296948 516284 296954
rect 516232 296890 516284 296896
rect 516140 296880 516192 296886
rect 516140 296822 516192 296828
rect 516152 295322 516180 296822
rect 516140 295316 516192 295322
rect 516140 295258 516192 295264
rect 516152 295089 516180 295258
rect 516244 295186 516272 296890
rect 516336 295254 516364 297502
rect 516416 297016 516468 297022
rect 516416 296958 516468 296964
rect 516324 295248 516376 295254
rect 516324 295190 516376 295196
rect 516232 295180 516284 295186
rect 516232 295122 516284 295128
rect 516138 295080 516194 295089
rect 516138 295015 516194 295024
rect 516244 294545 516272 295122
rect 516230 294536 516286 294545
rect 516230 294471 516286 294480
rect 516336 294001 516364 295190
rect 516322 293992 516378 294001
rect 516232 293956 516284 293962
rect 516322 293927 516378 293936
rect 516232 293898 516284 293904
rect 516140 293888 516192 293894
rect 516244 293865 516272 293898
rect 516140 293830 516192 293836
rect 516230 293856 516286 293865
rect 516152 293457 516180 293830
rect 516230 293791 516286 293800
rect 516138 293448 516194 293457
rect 516138 293383 516194 293392
rect 516244 292913 516272 293791
rect 516230 292904 516286 292913
rect 516230 292839 516286 292848
rect 516324 292528 516376 292534
rect 516324 292470 516376 292476
rect 516140 292460 516192 292466
rect 516140 292402 516192 292408
rect 516152 292369 516180 292402
rect 516232 292392 516284 292398
rect 516138 292360 516194 292369
rect 516232 292334 516284 292340
rect 516138 292295 516194 292304
rect 516244 291281 516272 292334
rect 516336 291825 516364 292470
rect 516322 291816 516378 291825
rect 516322 291751 516378 291760
rect 516230 291272 516286 291281
rect 516230 291207 516286 291216
rect 516324 291168 516376 291174
rect 516324 291110 516376 291116
rect 516232 291100 516284 291106
rect 516232 291042 516284 291048
rect 516244 290737 516272 291042
rect 516230 290728 516286 290737
rect 516230 290663 516286 290672
rect 516336 290193 516364 291110
rect 516322 290184 516378 290193
rect 516322 290119 516378 290128
rect 516324 289808 516376 289814
rect 516324 289750 516376 289756
rect 516232 289740 516284 289746
rect 516232 289682 516284 289688
rect 516140 289672 516192 289678
rect 516138 289640 516140 289649
rect 516192 289640 516194 289649
rect 516138 289575 516194 289584
rect 516244 289105 516272 289682
rect 516230 289096 516286 289105
rect 516230 289031 516286 289040
rect 516336 288561 516364 289750
rect 516322 288552 516378 288561
rect 516322 288487 516378 288496
rect 516428 285433 516456 296958
rect 516520 289814 516548 298318
rect 516612 292534 516640 298726
rect 516692 298444 516744 298450
rect 516692 298386 516744 298392
rect 516600 292528 516652 292534
rect 516600 292470 516652 292476
rect 516704 291106 516732 298386
rect 516796 291174 516824 298794
rect 516980 297809 517008 306346
rect 516966 297800 517022 297809
rect 516966 297735 517022 297744
rect 516784 291168 516836 291174
rect 516784 291110 516836 291116
rect 516692 291100 516744 291106
rect 516692 291042 516744 291048
rect 516508 289808 516560 289814
rect 516508 289750 516560 289756
rect 516414 285424 516470 285433
rect 516414 285359 516470 285368
rect 516782 284880 516838 284889
rect 516782 284815 516838 284824
rect 516506 284336 516562 284345
rect 516506 284271 516562 284280
rect 516414 283792 516470 283801
rect 516414 283727 516470 283736
rect 516322 282704 516378 282713
rect 516322 282639 516378 282648
rect 516138 281616 516194 281625
rect 516138 281551 516140 281560
rect 516192 281551 516194 281560
rect 516140 281522 516192 281528
rect 516230 281072 516286 281081
rect 516230 281007 516286 281016
rect 516138 280528 516194 280537
rect 516138 280463 516140 280472
rect 516192 280463 516194 280472
rect 516140 280434 516192 280440
rect 516244 280226 516272 281007
rect 516232 280220 516284 280226
rect 516232 280162 516284 280168
rect 516230 279984 516286 279993
rect 516230 279919 516286 279928
rect 516138 279440 516194 279449
rect 516138 279375 516194 279384
rect 516152 278866 516180 279375
rect 516140 278860 516192 278866
rect 516140 278802 516192 278808
rect 516244 278798 516272 279919
rect 516232 278792 516284 278798
rect 516232 278734 516284 278740
rect 516140 278724 516192 278730
rect 516140 278666 516192 278672
rect 516152 276962 516180 278666
rect 516336 278610 516364 282639
rect 516428 278730 516456 283727
rect 516416 278724 516468 278730
rect 516416 278666 516468 278672
rect 516244 278582 516364 278610
rect 516140 276956 516192 276962
rect 516140 276898 516192 276904
rect 516138 276856 516194 276865
rect 516138 276791 516140 276800
rect 516192 276791 516194 276800
rect 516140 276762 516192 276768
rect 516140 275256 516192 275262
rect 516138 275224 516140 275233
rect 516192 275224 516194 275233
rect 516138 275159 516194 275168
rect 516140 274712 516192 274718
rect 516138 274680 516140 274689
rect 516192 274680 516194 274689
rect 516138 274615 516194 274624
rect 516140 273216 516192 273222
rect 516140 273158 516192 273164
rect 516152 273057 516180 273158
rect 516138 273048 516194 273057
rect 516138 272983 516194 272992
rect 516138 271960 516194 271969
rect 516138 271895 516140 271904
rect 516192 271895 516194 271904
rect 516140 271866 516192 271872
rect 516138 271416 516194 271425
rect 516138 271351 516194 271360
rect 516152 271250 516180 271351
rect 516140 271244 516192 271250
rect 516140 271186 516192 271192
rect 516140 270224 516192 270230
rect 516140 270166 516192 270172
rect 516152 269793 516180 270166
rect 516138 269784 516194 269793
rect 516138 269719 516194 269728
rect 516138 269240 516194 269249
rect 516138 269175 516194 269184
rect 516152 269142 516180 269175
rect 516140 269136 516192 269142
rect 516140 269078 516192 269084
rect 516138 268696 516194 268705
rect 516138 268631 516140 268640
rect 516192 268631 516194 268640
rect 516140 268602 516192 268608
rect 516244 267714 516272 278582
rect 516414 278352 516470 278361
rect 516414 278287 516470 278296
rect 516428 277438 516456 278287
rect 516416 277432 516468 277438
rect 516322 277400 516378 277409
rect 516416 277374 516468 277380
rect 516322 277335 516378 277344
rect 516336 276078 516364 277335
rect 516416 276956 516468 276962
rect 516416 276898 516468 276904
rect 516324 276072 516376 276078
rect 516324 276014 516376 276020
rect 516322 275768 516378 275777
rect 516322 275703 516378 275712
rect 516336 275194 516364 275703
rect 516324 275188 516376 275194
rect 516324 275130 516376 275136
rect 516324 272536 516376 272542
rect 516322 272504 516324 272513
rect 516376 272504 516378 272513
rect 516322 272439 516378 272448
rect 516324 271176 516376 271182
rect 516324 271118 516376 271124
rect 516336 270881 516364 271118
rect 516322 270872 516378 270881
rect 516322 270807 516378 270816
rect 516322 270328 516378 270337
rect 516322 270263 516378 270272
rect 516336 269550 516364 270263
rect 516324 269544 516376 269550
rect 516324 269486 516376 269492
rect 516428 268530 516456 276898
rect 516520 268598 516548 284271
rect 516598 283248 516654 283257
rect 516598 283183 516654 283192
rect 516508 268592 516560 268598
rect 516508 268534 516560 268540
rect 516416 268524 516468 268530
rect 516416 268466 516468 268472
rect 516612 268462 516640 283183
rect 516690 277944 516746 277953
rect 516690 277879 516692 277888
rect 516744 277879 516746 277888
rect 516692 277850 516744 277856
rect 516692 276344 516744 276350
rect 516690 276312 516692 276321
rect 516744 276312 516746 276321
rect 516690 276247 516746 276256
rect 516690 274136 516746 274145
rect 516690 274071 516692 274080
rect 516744 274071 516746 274080
rect 516692 274042 516744 274048
rect 516600 268456 516652 268462
rect 516600 268398 516652 268404
rect 516796 268394 516824 284815
rect 516980 277394 517008 297735
rect 517152 297356 517204 297362
rect 517152 297298 517204 297304
rect 517058 296712 517114 296721
rect 517058 296647 517114 296656
rect 516888 277366 517008 277394
rect 516784 268388 516836 268394
rect 516784 268330 516836 268336
rect 516232 267708 516284 267714
rect 516232 267650 516284 267656
rect 516232 234592 516284 234598
rect 516232 234534 516284 234540
rect 516244 233306 516272 234534
rect 516232 233300 516284 233306
rect 516232 233242 516284 233248
rect 516600 233300 516652 233306
rect 516600 233242 516652 233248
rect 516416 233232 516468 233238
rect 516416 233174 516468 233180
rect 516428 231878 516456 233174
rect 516416 231872 516468 231878
rect 516416 231814 516468 231820
rect 516232 226840 516284 226846
rect 516232 226782 516284 226788
rect 516244 226370 516272 226782
rect 516232 226364 516284 226370
rect 516232 226306 516284 226312
rect 516140 226296 516192 226302
rect 516140 226238 516192 226244
rect 516152 225457 516180 226238
rect 516138 225448 516194 225457
rect 516138 225383 516194 225392
rect 516140 224936 516192 224942
rect 516140 224878 516192 224884
rect 516152 224369 516180 224878
rect 516138 224360 516194 224369
rect 516138 224295 516194 224304
rect 516140 222148 516192 222154
rect 516140 222090 516192 222096
rect 516152 222057 516180 222090
rect 516138 222048 516194 222057
rect 516138 221983 516194 221992
rect 516138 220824 516194 220833
rect 516138 220759 516140 220768
rect 516192 220759 516194 220768
rect 516140 220730 516192 220736
rect 516140 219972 516192 219978
rect 516140 219914 516192 219920
rect 516152 219745 516180 219914
rect 516138 219736 516194 219745
rect 516138 219671 516194 219680
rect 516140 219360 516192 219366
rect 516140 219302 516192 219308
rect 516152 218521 516180 219302
rect 516138 218512 516194 218521
rect 516138 218447 516194 218456
rect 516428 217433 516456 231814
rect 516508 226364 516560 226370
rect 516508 226306 516560 226312
rect 516414 217424 516470 217433
rect 516414 217359 516470 217368
rect 516140 216640 516192 216646
rect 516140 216582 516192 216588
rect 516152 216209 516180 216582
rect 516138 216200 516194 216209
rect 516138 216135 516194 216144
rect 516520 215121 516548 226306
rect 516612 223145 516640 233242
rect 516598 223136 516654 223145
rect 516598 223071 516654 223080
rect 516506 215112 516562 215121
rect 516506 215047 516562 215056
rect 516232 213920 516284 213926
rect 516230 213888 516232 213897
rect 516284 213888 516286 213897
rect 516140 213852 516192 213858
rect 516230 213823 516286 213832
rect 516140 213794 516192 213800
rect 516152 212809 516180 213794
rect 516138 212800 516194 212809
rect 516138 212735 516194 212744
rect 516140 211948 516192 211954
rect 516140 211890 516192 211896
rect 516152 211585 516180 211890
rect 516138 211576 516194 211585
rect 516138 211511 516194 211520
rect 516140 209568 516192 209574
rect 516140 209510 516192 209516
rect 516152 209273 516180 209510
rect 516138 209264 516194 209273
rect 516138 209199 516194 209208
rect 516138 206952 516194 206961
rect 516138 206887 516140 206896
rect 516192 206887 516194 206896
rect 516140 206858 516192 206864
rect 515404 206848 515456 206854
rect 515404 206790 515456 206796
rect 516140 205896 516192 205902
rect 516138 205864 516140 205873
rect 516192 205864 516194 205873
rect 516138 205799 516194 205808
rect 516140 204944 516192 204950
rect 516140 204886 516192 204892
rect 516152 204649 516180 204886
rect 516138 204640 516194 204649
rect 516138 204575 516194 204584
rect 516140 204264 516192 204270
rect 516140 204206 516192 204212
rect 516152 203561 516180 204206
rect 516138 203552 516194 203561
rect 516138 203487 516194 203496
rect 516140 202836 516192 202842
rect 516140 202778 516192 202784
rect 516152 202337 516180 202778
rect 516138 202328 516194 202337
rect 516138 202263 516194 202272
rect 516244 200114 516272 213823
rect 516416 211132 516468 211138
rect 516416 211074 516468 211080
rect 516428 210497 516456 211074
rect 516414 210488 516470 210497
rect 516414 210423 516470 210432
rect 516428 209774 516456 210423
rect 516428 209746 516548 209774
rect 516324 204944 516376 204950
rect 516324 204886 516376 204892
rect 516152 200086 516272 200114
rect 514944 197328 514996 197334
rect 514944 197270 514996 197276
rect 516152 196654 516180 200086
rect 516336 197198 516364 204886
rect 516520 197266 516548 209746
rect 516508 197260 516560 197266
rect 516508 197202 516560 197208
rect 516324 197192 516376 197198
rect 516324 197134 516376 197140
rect 516140 196648 516192 196654
rect 516140 196590 516192 196596
rect 508872 194404 508924 194410
rect 508872 194346 508924 194352
rect 514852 194404 514904 194410
rect 514852 194346 514904 194352
rect 513380 156256 513432 156262
rect 513380 156198 513432 156204
rect 507768 155304 507820 155310
rect 507768 155246 507820 155252
rect 513196 154012 513248 154018
rect 513196 153954 513248 153960
rect 513104 151972 513156 151978
rect 513104 151914 513156 151920
rect 513116 142746 513144 151914
rect 513208 148866 513236 153954
rect 513288 153196 513340 153202
rect 513288 153138 513340 153144
rect 513300 149025 513328 153138
rect 513392 152969 513420 156198
rect 515036 156188 515088 156194
rect 515036 156130 515088 156136
rect 513930 156088 513986 156097
rect 513930 156023 513986 156032
rect 513656 154148 513708 154154
rect 513656 154090 513708 154096
rect 513562 153912 513618 153921
rect 513562 153847 513618 153856
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 513378 152960 513434 152969
rect 513378 152895 513434 152904
rect 513380 152788 513432 152794
rect 513380 152730 513432 152736
rect 513392 149705 513420 152730
rect 513378 149696 513434 149705
rect 513378 149631 513434 149640
rect 513286 149016 513342 149025
rect 513286 148951 513342 148960
rect 513208 148838 513420 148866
rect 513392 148458 513420 148838
rect 513484 148617 513512 153070
rect 513576 151745 513604 153847
rect 513562 151736 513618 151745
rect 513562 151671 513618 151680
rect 513564 151632 513616 151638
rect 513564 151574 513616 151580
rect 513470 148608 513526 148617
rect 513470 148543 513526 148552
rect 513392 148430 513512 148458
rect 513380 147144 513432 147150
rect 513380 147086 513432 147092
rect 513286 142760 513342 142769
rect 513116 142718 513286 142746
rect 513286 142695 513342 142704
rect 503076 135312 503128 135318
rect 503076 135254 503128 135260
rect 503088 124098 503116 135254
rect 513392 134065 513420 147086
rect 513378 134056 513434 134065
rect 513378 133991 513434 134000
rect 503168 133952 503220 133958
rect 503168 133894 503220 133900
rect 503076 124092 503128 124098
rect 503076 124034 503128 124040
rect 503180 124030 503208 133894
rect 503260 132524 503312 132530
rect 503260 132466 503312 132472
rect 503168 124024 503220 124030
rect 503168 123966 503220 123972
rect 503272 123894 503300 132466
rect 513484 132433 513512 148430
rect 513576 147150 513604 151574
rect 513668 151337 513696 154090
rect 513748 154080 513800 154086
rect 513748 154022 513800 154028
rect 513654 151328 513710 151337
rect 513654 151263 513710 151272
rect 513760 150249 513788 154022
rect 513840 153672 513892 153678
rect 513840 153614 513892 153620
rect 513852 152425 513880 153614
rect 513838 152416 513894 152425
rect 513838 152351 513894 152360
rect 513944 152266 513972 156023
rect 514024 155304 514076 155310
rect 514024 155246 514076 155252
rect 513852 152238 513972 152266
rect 513746 150240 513802 150249
rect 513746 150175 513802 150184
rect 513564 147144 513616 147150
rect 513564 147086 513616 147092
rect 513656 147076 513708 147082
rect 513656 147018 513708 147024
rect 513564 147008 513616 147014
rect 513564 146950 513616 146956
rect 513470 132424 513526 132433
rect 513470 132359 513526 132368
rect 513576 131481 513604 146950
rect 513668 133657 513696 147018
rect 513748 146940 513800 146946
rect 513748 146882 513800 146888
rect 513654 133648 513710 133657
rect 513654 133583 513710 133592
rect 513760 133113 513788 146882
rect 513852 136649 513880 152238
rect 513932 152176 513984 152182
rect 513932 152118 513984 152124
rect 513944 137329 513972 152118
rect 513930 137320 513986 137329
rect 513930 137255 513986 137264
rect 513838 136640 513894 136649
rect 513838 136575 513894 136584
rect 513746 133104 513802 133113
rect 513746 133039 513802 133048
rect 513562 131472 513618 131481
rect 513562 131407 513618 131416
rect 513286 129160 513342 129169
rect 513286 129095 513342 129104
rect 503628 129056 503680 129062
rect 503628 128998 503680 129004
rect 503640 123962 503668 128998
rect 504272 127696 504324 127702
rect 504272 127638 504324 127644
rect 503628 123956 503680 123962
rect 503628 123898 503680 123904
rect 503260 123888 503312 123894
rect 503260 123830 503312 123836
rect 504284 123758 504312 127638
rect 504364 127628 504416 127634
rect 504364 127570 504416 127576
rect 504376 123826 504404 127570
rect 513196 125248 513248 125254
rect 513196 125190 513248 125196
rect 513208 124386 513236 125190
rect 513300 125050 513328 129095
rect 513470 128616 513526 128625
rect 513470 128551 513526 128560
rect 513378 125352 513434 125361
rect 513378 125287 513434 125296
rect 513392 125186 513420 125287
rect 513380 125180 513432 125186
rect 513380 125122 513432 125128
rect 513288 125044 513340 125050
rect 513288 124986 513340 124992
rect 513380 125044 513432 125050
rect 513380 124986 513432 124992
rect 513392 124953 513420 124986
rect 513378 124944 513434 124953
rect 513484 124914 513512 128551
rect 513838 128072 513894 128081
rect 513838 128007 513894 128016
rect 513746 127528 513802 127537
rect 513746 127463 513802 127472
rect 513654 125896 513710 125905
rect 513654 125831 513710 125840
rect 513562 125352 513618 125361
rect 513562 125287 513618 125296
rect 513378 124879 513434 124888
rect 513472 124908 513524 124914
rect 513472 124850 513524 124856
rect 513286 124400 513342 124409
rect 513208 124358 513286 124386
rect 513286 124335 513342 124344
rect 504364 123820 504416 123826
rect 504364 123762 504416 123768
rect 504272 123752 504324 123758
rect 504272 123694 504324 123700
rect 504928 122738 504956 124100
rect 506860 122738 506888 124100
rect 504916 122732 504968 122738
rect 504916 122674 504968 122680
rect 506848 122732 506900 122738
rect 506848 122674 506900 122680
rect 508884 122670 508912 124100
rect 510908 122874 510936 124100
rect 510896 122868 510948 122874
rect 510896 122810 510948 122816
rect 512932 122806 512960 124100
rect 513576 123962 513604 125287
rect 513564 123956 513616 123962
rect 513564 123898 513616 123904
rect 513668 123826 513696 125831
rect 513760 124030 513788 127463
rect 513852 124098 513880 128007
rect 513930 127120 513986 127129
rect 513930 127055 513986 127064
rect 513840 124092 513892 124098
rect 513840 124034 513892 124040
rect 513748 124024 513800 124030
rect 513748 123966 513800 123972
rect 513944 123894 513972 127055
rect 513932 123888 513984 123894
rect 513932 123830 513984 123836
rect 513656 123820 513708 123826
rect 513656 123762 513708 123768
rect 512920 122800 512972 122806
rect 512920 122742 512972 122748
rect 514036 122738 514064 155246
rect 514116 154216 514168 154222
rect 514116 154158 514168 154164
rect 514128 151774 514156 154158
rect 514392 153808 514444 153814
rect 514392 153750 514444 153756
rect 514208 153536 514260 153542
rect 514208 153478 514260 153484
rect 514116 151768 514168 151774
rect 514116 151710 514168 151716
rect 514220 151706 514248 153478
rect 514300 153468 514352 153474
rect 514300 153410 514352 153416
rect 514208 151700 514260 151706
rect 514208 151642 514260 151648
rect 514312 151586 514340 153410
rect 514404 152017 514432 153750
rect 514576 153740 514628 153746
rect 514576 153682 514628 153688
rect 514484 153604 514536 153610
rect 514484 153546 514536 153552
rect 514390 152008 514446 152017
rect 514390 151943 514446 151952
rect 514390 151872 514446 151881
rect 514390 151807 514446 151816
rect 514404 151706 514432 151807
rect 514392 151700 514444 151706
rect 514392 151642 514444 151648
rect 514312 151558 514432 151586
rect 514300 151496 514352 151502
rect 514206 151464 514262 151473
rect 514300 151438 514352 151444
rect 514206 151399 514262 151408
rect 514114 151328 514170 151337
rect 514114 151263 514170 151272
rect 514128 131753 514156 151263
rect 514220 135425 514248 151399
rect 514312 150793 514340 151438
rect 514298 150784 514354 150793
rect 514298 150719 514354 150728
rect 514300 150680 514352 150686
rect 514300 150622 514352 150628
rect 514312 146169 514340 150622
rect 514404 147014 514432 151558
rect 514496 147082 514524 153546
rect 514484 147076 514536 147082
rect 514484 147018 514536 147024
rect 514392 147008 514444 147014
rect 514392 146950 514444 146956
rect 514588 146946 514616 153682
rect 514760 153400 514812 153406
rect 514760 153342 514812 153348
rect 514668 153332 514720 153338
rect 514668 153274 514720 153280
rect 514576 146940 514628 146946
rect 514576 146882 514628 146888
rect 514298 146160 514354 146169
rect 514298 146095 514354 146104
rect 514680 142154 514708 153274
rect 514312 142126 514708 142154
rect 514312 141409 514340 142126
rect 514298 141400 514354 141409
rect 514298 141335 514354 141344
rect 514206 135416 514262 135425
rect 514206 135351 514262 135360
rect 514772 134337 514800 153342
rect 514944 152108 514996 152114
rect 514944 152050 514996 152056
rect 514852 152040 514904 152046
rect 514852 151982 514904 151988
rect 514864 134881 514892 151982
rect 514956 135969 514984 152050
rect 515048 140321 515076 156130
rect 515128 156120 515180 156126
rect 515128 156062 515180 156068
rect 515140 140865 515168 156062
rect 515312 156052 515364 156058
rect 515312 155994 515364 156000
rect 515220 154624 515272 154630
rect 515220 154566 515272 154572
rect 515232 141953 515260 154566
rect 515218 141944 515274 141953
rect 515218 141879 515274 141888
rect 515126 140856 515182 140865
rect 515126 140791 515182 140800
rect 515034 140312 515090 140321
rect 515034 140247 515090 140256
rect 515324 139777 515352 155994
rect 516600 155236 516652 155242
rect 516600 155178 516652 155184
rect 515404 153876 515456 153882
rect 515404 153818 515456 153824
rect 515416 144906 515444 153818
rect 515588 153264 515640 153270
rect 515588 153206 515640 153212
rect 515496 151904 515548 151910
rect 515496 151846 515548 151852
rect 515404 144900 515456 144906
rect 515404 144842 515456 144848
rect 515310 139768 515366 139777
rect 515310 139703 515366 139712
rect 515508 139233 515536 151846
rect 515600 143041 515628 153206
rect 516232 153128 516284 153134
rect 516232 153070 516284 153076
rect 516140 153060 516192 153066
rect 516140 153002 516192 153008
rect 516152 152697 516180 153002
rect 516138 152688 516194 152697
rect 516138 152623 516194 152632
rect 516140 152584 516192 152590
rect 516140 152526 516192 152532
rect 516152 145625 516180 152526
rect 516244 152153 516272 153070
rect 516508 152856 516560 152862
rect 516508 152798 516560 152804
rect 516324 152720 516376 152726
rect 516324 152662 516376 152668
rect 516230 152144 516286 152153
rect 516230 152079 516286 152088
rect 516336 151994 516364 152662
rect 516416 152516 516468 152522
rect 516416 152458 516468 152464
rect 516244 151966 516364 151994
rect 516244 147257 516272 151966
rect 516324 151904 516376 151910
rect 516324 151846 516376 151852
rect 516336 147801 516364 151846
rect 516322 147792 516378 147801
rect 516322 147727 516378 147736
rect 516230 147248 516286 147257
rect 516230 147183 516286 147192
rect 516138 145616 516194 145625
rect 516138 145551 516194 145560
rect 516428 145081 516456 152458
rect 516520 151978 516548 152798
rect 516508 151972 516560 151978
rect 516508 151914 516560 151920
rect 516508 151836 516560 151842
rect 516508 151778 516560 151784
rect 516414 145072 516470 145081
rect 516414 145007 516470 145016
rect 516140 144900 516192 144906
rect 516140 144842 516192 144848
rect 515586 143032 515642 143041
rect 515586 142967 515642 142976
rect 515494 139224 515550 139233
rect 515494 139159 515550 139168
rect 516152 137601 516180 144842
rect 516520 143585 516548 151778
rect 516612 144537 516640 155178
rect 516784 153944 516836 153950
rect 516784 153886 516836 153892
rect 516692 152924 516744 152930
rect 516692 152866 516744 152872
rect 516704 146713 516732 152866
rect 516690 146704 516746 146713
rect 516690 146639 516746 146648
rect 516598 144528 516654 144537
rect 516598 144463 516654 144472
rect 516796 144129 516824 153886
rect 516888 153785 516916 277366
rect 517072 217394 517100 296647
rect 517164 282169 517192 297298
rect 517256 296614 517284 439991
rect 517348 297265 517376 441079
rect 517426 417480 517482 417489
rect 517532 417466 517560 495450
rect 517610 484664 517666 484673
rect 517610 484599 517666 484608
rect 517482 417438 517560 417466
rect 517426 417415 517482 417424
rect 517426 352200 517482 352209
rect 517532 352186 517560 417438
rect 517624 412185 517652 484599
rect 517704 439136 517756 439142
rect 517704 439078 517756 439084
rect 517716 417382 517744 439078
rect 518176 425746 518204 514014
rect 518900 510672 518952 510678
rect 518900 510614 518952 510620
rect 518256 501424 518308 501430
rect 518256 501366 518308 501372
rect 518164 425740 518216 425746
rect 518164 425682 518216 425688
rect 517796 424584 517848 424590
rect 517796 424526 517848 424532
rect 517704 417376 517756 417382
rect 517704 417318 517756 417324
rect 517610 412176 517666 412185
rect 517610 412111 517666 412120
rect 517808 368422 517836 424526
rect 517888 421932 517940 421938
rect 517888 421874 517940 421880
rect 517900 389230 517928 421874
rect 518268 420238 518296 501366
rect 518912 424454 518940 510614
rect 519004 500818 519032 563246
rect 519084 562556 519136 562562
rect 519084 562498 519136 562504
rect 518992 500812 519044 500818
rect 518992 500754 519044 500760
rect 518900 424448 518952 424454
rect 518900 424390 518952 424396
rect 518256 420232 518308 420238
rect 518256 420174 518308 420180
rect 519004 420034 519032 500754
rect 519096 498506 519124 562498
rect 519176 557796 519228 557802
rect 519176 557738 519228 557744
rect 519084 498500 519136 498506
rect 519084 498442 519136 498448
rect 518072 420028 518124 420034
rect 518072 419970 518124 419976
rect 518992 420028 519044 420034
rect 518992 419970 519044 419976
rect 517980 417444 518032 417450
rect 517980 417386 518032 417392
rect 517888 389224 517940 389230
rect 517888 389166 517940 389172
rect 517796 368416 517848 368422
rect 517796 368358 517848 368364
rect 517900 362710 517928 389166
rect 517888 362704 517940 362710
rect 517888 362646 517940 362652
rect 517992 354674 518020 417386
rect 518084 357406 518112 419970
rect 518900 419824 518952 419830
rect 518900 419766 518952 419772
rect 518256 360868 518308 360874
rect 518256 360810 518308 360816
rect 518072 357400 518124 357406
rect 518072 357342 518124 357348
rect 517624 354646 518020 354674
rect 517624 353297 517652 354646
rect 517610 353288 517666 353297
rect 517610 353223 517666 353232
rect 517482 352158 517560 352186
rect 517426 352135 517482 352144
rect 517334 297256 517390 297265
rect 517334 297191 517390 297200
rect 517244 296608 517296 296614
rect 517244 296550 517296 296556
rect 517256 296002 517284 296550
rect 517244 295996 517296 296002
rect 517244 295938 517296 295944
rect 517150 282160 517206 282169
rect 517150 282095 517206 282104
rect 517060 217388 517112 217394
rect 517060 217330 517112 217336
rect 517348 207074 517376 297191
rect 517426 273592 517482 273601
rect 517532 273578 517560 352158
rect 517624 274106 517652 353223
rect 517704 349852 517756 349858
rect 517704 349794 517756 349800
rect 517716 287054 517744 349794
rect 518164 299668 518216 299674
rect 518164 299610 518216 299616
rect 517716 287026 517928 287054
rect 517796 279472 517848 279478
rect 517796 279414 517848 279420
rect 517808 278905 517836 279414
rect 517794 278896 517850 278905
rect 517794 278831 517850 278840
rect 517612 274100 517664 274106
rect 517612 274042 517664 274048
rect 517482 273550 517560 273578
rect 517426 273527 517482 273536
rect 517532 273290 517560 273550
rect 517520 273284 517572 273290
rect 517520 273226 517572 273232
rect 517808 243574 517836 278831
rect 517900 272542 517928 287026
rect 518072 276344 518124 276350
rect 518072 276286 518124 276292
rect 517888 272536 517940 272542
rect 517888 272478 517940 272484
rect 517796 243568 517848 243574
rect 517796 243510 517848 243516
rect 517900 239426 517928 272478
rect 517980 243568 518032 243574
rect 517980 243510 518032 243516
rect 517888 239420 517940 239426
rect 517888 239362 517940 239368
rect 517900 238754 517928 239362
rect 517808 238726 517928 238754
rect 517704 228744 517756 228750
rect 517704 228686 517756 228692
rect 517716 228478 517744 228686
rect 517704 228472 517756 228478
rect 517704 228414 517756 228420
rect 517716 209774 517744 228414
rect 517532 209746 517744 209774
rect 517426 208176 517482 208185
rect 517532 208162 517560 209746
rect 517482 208134 517560 208162
rect 517426 208111 517482 208120
rect 517348 207046 517560 207074
rect 517532 200114 517560 207046
rect 517808 205902 517836 238726
rect 517992 219978 518020 243510
rect 517980 219972 518032 219978
rect 517980 219914 518032 219920
rect 518084 213926 518112 276286
rect 518072 213920 518124 213926
rect 518072 213862 518124 213868
rect 517796 205896 517848 205902
rect 517796 205838 517848 205844
rect 517532 200086 517652 200114
rect 517426 196616 517482 196625
rect 517482 196574 517560 196602
rect 517426 196551 517482 196560
rect 516968 155984 517020 155990
rect 516968 155926 517020 155932
rect 516874 153776 516930 153785
rect 516874 153711 516930 153720
rect 516980 151842 517008 155926
rect 516968 151836 517020 151842
rect 516968 151778 517020 151784
rect 516782 144120 516838 144129
rect 516782 144055 516838 144064
rect 516506 143576 516562 143585
rect 516506 143511 516562 143520
rect 516506 138680 516562 138689
rect 516506 138615 516562 138624
rect 516230 138136 516286 138145
rect 516230 138071 516286 138080
rect 516138 137592 516194 137601
rect 516138 137527 516194 137536
rect 514942 135960 514998 135969
rect 514942 135895 514998 135904
rect 514850 134872 514906 134881
rect 514850 134807 514906 134816
rect 514758 134328 514814 134337
rect 514758 134263 514814 134272
rect 516244 132494 516272 138071
rect 516244 132466 516364 132494
rect 514114 131744 514170 131753
rect 514114 131679 514170 131688
rect 516138 130656 516194 130665
rect 516138 130591 516194 130600
rect 514114 126440 514170 126449
rect 514114 126375 514170 126384
rect 514128 123758 514156 126375
rect 516152 124982 516180 130591
rect 516230 130112 516286 130121
rect 516230 130047 516286 130056
rect 516140 124976 516192 124982
rect 516140 124918 516192 124924
rect 516244 124846 516272 130047
rect 516232 124840 516284 124846
rect 516232 124782 516284 124788
rect 516336 124778 516364 132466
rect 516324 124772 516376 124778
rect 516324 124714 516376 124720
rect 516520 124166 516548 138615
rect 517426 124264 517482 124273
rect 517532 124250 517560 196574
rect 517624 153241 517652 200086
rect 517610 153232 517666 153241
rect 517610 153167 517666 153176
rect 518176 139398 518204 299610
rect 518268 277914 518296 360810
rect 518912 359174 518940 419766
rect 518992 418600 519044 418606
rect 518992 418542 519044 418548
rect 518900 359168 518952 359174
rect 518900 359110 518952 359116
rect 519004 355638 519032 418542
rect 519096 418538 519124 498442
rect 519188 491230 519216 557738
rect 519280 516118 519308 564470
rect 519268 516112 519320 516118
rect 519268 516054 519320 516060
rect 519372 508842 519400 567258
rect 520280 563780 520332 563786
rect 520280 563722 520332 563728
rect 519360 508836 519412 508842
rect 519360 508778 519412 508784
rect 519372 507890 519400 508778
rect 519360 507884 519412 507890
rect 519360 507826 519412 507832
rect 520292 501430 520320 563722
rect 520384 512786 520412 568890
rect 521752 567384 521804 567390
rect 521752 567326 521804 567332
rect 520464 566092 520516 566098
rect 520464 566034 520516 566040
rect 520476 517546 520504 566034
rect 520556 564732 520608 564738
rect 520556 564674 520608 564680
rect 520568 536110 520596 564674
rect 521660 556300 521712 556306
rect 521660 556242 521712 556248
rect 520556 536104 520608 536110
rect 520556 536046 520608 536052
rect 520464 517540 520516 517546
rect 520464 517482 520516 517488
rect 520372 512780 520424 512786
rect 520372 512722 520424 512728
rect 520372 505436 520424 505442
rect 520372 505378 520424 505384
rect 520280 501424 520332 501430
rect 520280 501366 520332 501372
rect 519176 491224 519228 491230
rect 519176 491166 519228 491172
rect 519176 423632 519228 423638
rect 519176 423574 519228 423580
rect 519188 422550 519216 423574
rect 519176 422544 519228 422550
rect 519176 422486 519228 422492
rect 519084 418532 519136 418538
rect 519084 418474 519136 418480
rect 519096 376038 519124 418474
rect 519084 376032 519136 376038
rect 519084 375974 519136 375980
rect 518992 355632 519044 355638
rect 518992 355574 519044 355580
rect 519004 287054 519032 355574
rect 519096 354550 519124 375974
rect 519188 371754 519216 422486
rect 520384 421598 520412 505378
rect 520568 505102 520596 536046
rect 520648 507884 520700 507890
rect 520648 507826 520700 507832
rect 520556 505096 520608 505102
rect 520556 505038 520608 505044
rect 520464 424448 520516 424454
rect 520464 424390 520516 424396
rect 520372 421592 520424 421598
rect 520372 421534 520424 421540
rect 520384 420986 520412 421534
rect 520372 420980 520424 420986
rect 520372 420922 520424 420928
rect 520280 420232 520332 420238
rect 520280 420174 520332 420180
rect 519544 414724 519596 414730
rect 519544 414666 519596 414672
rect 519176 371748 519228 371754
rect 519176 371690 519228 371696
rect 519176 359168 519228 359174
rect 519176 359110 519228 359116
rect 519084 354544 519136 354550
rect 519084 354486 519136 354492
rect 519004 287026 519124 287054
rect 518900 280492 518952 280498
rect 518900 280434 518952 280440
rect 518256 277908 518308 277914
rect 518256 277850 518308 277856
rect 518268 277506 518296 277850
rect 518256 277500 518308 277506
rect 518256 277442 518308 277448
rect 518348 274712 518400 274718
rect 518348 274654 518400 274660
rect 518256 273284 518308 273290
rect 518256 273226 518308 273232
rect 518268 228750 518296 273226
rect 518256 228744 518308 228750
rect 518256 228686 518308 228692
rect 518360 211138 518388 274654
rect 518912 234598 518940 280434
rect 519096 275262 519124 287026
rect 519188 276826 519216 359110
rect 519556 346322 519584 414666
rect 520292 357950 520320 420174
rect 520372 412548 520424 412554
rect 520372 412490 520424 412496
rect 520280 357944 520332 357950
rect 520280 357886 520332 357892
rect 519544 346316 519596 346322
rect 519544 346258 519596 346264
rect 519636 344344 519688 344350
rect 519636 344286 519688 344292
rect 519544 301028 519596 301034
rect 519544 300970 519596 300976
rect 519268 277500 519320 277506
rect 519268 277442 519320 277448
rect 519176 276820 519228 276826
rect 519176 276762 519228 276768
rect 519188 276146 519216 276762
rect 519176 276140 519228 276146
rect 519176 276082 519228 276088
rect 519084 275256 519136 275262
rect 519084 275198 519136 275204
rect 519096 236706 519124 275198
rect 519176 274100 519228 274106
rect 519176 274042 519228 274048
rect 519188 240786 519216 274042
rect 519176 240780 519228 240786
rect 519176 240722 519228 240728
rect 519084 236700 519136 236706
rect 519084 236642 519136 236648
rect 518900 234592 518952 234598
rect 518900 234534 518952 234540
rect 518900 217388 518952 217394
rect 518900 217330 518952 217336
rect 518348 211132 518400 211138
rect 518348 211074 518400 211080
rect 518912 153066 518940 217330
rect 519096 211954 519124 236642
rect 519084 211948 519136 211954
rect 519084 211890 519136 211896
rect 519188 209574 519216 240722
rect 519280 233238 519308 277442
rect 519268 233232 519320 233238
rect 519268 233174 519320 233180
rect 519556 219434 519584 300970
rect 519648 270230 519676 344286
rect 520292 276350 520320 357886
rect 520384 341766 520412 412490
rect 520476 367810 520504 424390
rect 520660 423638 520688 507826
rect 520924 486464 520976 486470
rect 520924 486406 520976 486412
rect 520648 423632 520700 423638
rect 520648 423574 520700 423580
rect 520648 421184 520700 421190
rect 520648 421126 520700 421132
rect 520556 415812 520608 415818
rect 520556 415754 520608 415760
rect 520568 373318 520596 415754
rect 520660 381546 520688 421126
rect 520936 413302 520964 486406
rect 521672 485790 521700 556242
rect 521764 509930 521792 567326
rect 521936 565888 521988 565894
rect 521936 565830 521988 565836
rect 521844 557660 521896 557666
rect 521844 557602 521896 557608
rect 521752 509924 521804 509930
rect 521752 509866 521804 509872
rect 521660 485784 521712 485790
rect 521660 485726 521712 485732
rect 521764 441614 521792 509866
rect 521856 489870 521884 557602
rect 521948 541686 521976 565830
rect 523040 557728 523092 557734
rect 523040 557670 523092 557676
rect 521936 541680 521988 541686
rect 521936 541622 521988 541628
rect 521948 507822 521976 541622
rect 521936 507816 521988 507822
rect 521936 507758 521988 507764
rect 522120 491224 522172 491230
rect 522120 491166 522172 491172
rect 521844 489864 521896 489870
rect 521844 489806 521896 489812
rect 521764 441586 522068 441614
rect 521660 434852 521712 434858
rect 521660 434794 521712 434800
rect 520924 413296 520976 413302
rect 520924 413238 520976 413244
rect 520648 381540 520700 381546
rect 520648 381482 520700 381488
rect 520556 373312 520608 373318
rect 520556 373254 520608 373260
rect 520464 367804 520516 367810
rect 520464 367746 520516 367752
rect 520568 348838 520596 373254
rect 520660 360738 520688 381482
rect 520648 360732 520700 360738
rect 520648 360674 520700 360680
rect 520556 348832 520608 348838
rect 520556 348774 520608 348780
rect 521016 347744 521068 347750
rect 521016 347686 521068 347692
rect 521028 347070 521056 347686
rect 521016 347064 521068 347070
rect 521016 347006 521068 347012
rect 520372 341760 520424 341766
rect 520372 341702 520424 341708
rect 520280 276344 520332 276350
rect 520280 276286 520332 276292
rect 519636 270224 519688 270230
rect 519636 270166 519688 270172
rect 520384 268666 520412 341702
rect 520924 302524 520976 302530
rect 520924 302466 520976 302472
rect 520464 276140 520516 276146
rect 520464 276082 520516 276088
rect 520372 268660 520424 268666
rect 520372 268602 520424 268608
rect 520384 258074 520412 268602
rect 520292 258046 520412 258074
rect 519544 219428 519596 219434
rect 519544 219370 519596 219376
rect 519176 209568 519228 209574
rect 519176 209510 519228 209516
rect 520292 198694 520320 258046
rect 520476 226846 520504 276082
rect 520556 275188 520608 275194
rect 520556 275130 520608 275136
rect 520568 229770 520596 275130
rect 520648 269544 520700 269550
rect 520648 269486 520700 269492
rect 520556 229764 520608 229770
rect 520556 229706 520608 229712
rect 520464 226840 520516 226846
rect 520464 226782 520516 226788
rect 520568 213858 520596 229706
rect 520556 213852 520608 213858
rect 520556 213794 520608 213800
rect 520660 201278 520688 269486
rect 520648 201272 520700 201278
rect 520648 201214 520700 201220
rect 520280 198688 520332 198694
rect 520280 198630 520332 198636
rect 520936 153202 520964 302466
rect 521028 271250 521056 347006
rect 521672 318102 521700 434794
rect 522040 424386 522068 441586
rect 522028 424380 522080 424386
rect 522028 424322 522080 424328
rect 521936 422340 521988 422346
rect 521936 422282 521988 422288
rect 521752 420980 521804 420986
rect 521752 420922 521804 420928
rect 521764 360874 521792 420922
rect 521844 412684 521896 412690
rect 521844 412626 521896 412632
rect 521752 360868 521804 360874
rect 521752 360810 521804 360816
rect 521856 344350 521884 412626
rect 521948 363662 521976 422282
rect 522040 377466 522068 424322
rect 522132 414730 522160 491166
rect 523052 488510 523080 557670
rect 523040 488504 523092 488510
rect 523040 488446 523092 488452
rect 524432 441590 524460 583714
rect 524604 568608 524656 568614
rect 524604 568550 524656 568556
rect 524512 556232 524564 556238
rect 524512 556174 524564 556180
rect 524524 486470 524552 556174
rect 524616 514078 524644 568550
rect 524696 559020 524748 559026
rect 524696 558962 524748 558968
rect 524708 522374 524736 558962
rect 525800 558952 525852 558958
rect 525800 558894 525852 558900
rect 525812 523734 525840 558894
rect 525800 523728 525852 523734
rect 525800 523670 525852 523676
rect 524696 522368 524748 522374
rect 524696 522310 524748 522316
rect 524604 514072 524656 514078
rect 524604 514014 524656 514020
rect 524708 492658 524736 522310
rect 525812 494018 525840 523670
rect 525800 494012 525852 494018
rect 525800 493954 525852 493960
rect 524696 492652 524748 492658
rect 524696 492594 524748 492600
rect 524512 486464 524564 486470
rect 524512 486406 524564 486412
rect 524420 441584 524472 441590
rect 524420 441526 524472 441532
rect 524420 437572 524472 437578
rect 524420 437514 524472 437520
rect 523040 436280 523092 436286
rect 523040 436222 523092 436228
rect 522120 414724 522172 414730
rect 522120 414666 522172 414672
rect 522028 377460 522080 377466
rect 522028 377402 522080 377408
rect 521936 363656 521988 363662
rect 521936 363598 521988 363604
rect 521844 344344 521896 344350
rect 521844 344286 521896 344292
rect 521660 318096 521712 318102
rect 521660 318038 521712 318044
rect 521672 292398 521700 318038
rect 521660 292392 521712 292398
rect 521660 292334 521712 292340
rect 521660 280220 521712 280226
rect 521660 280162 521712 280168
rect 521016 271244 521068 271250
rect 521016 271186 521068 271192
rect 521672 224942 521700 280162
rect 521948 279478 521976 363598
rect 522028 346316 522080 346322
rect 522028 346258 522080 346264
rect 521936 279472 521988 279478
rect 521936 279414 521988 279420
rect 521752 277432 521804 277438
rect 521752 277374 521804 277380
rect 521764 235278 521792 277374
rect 521936 276072 521988 276078
rect 521936 276014 521988 276020
rect 521844 271176 521896 271182
rect 521844 271118 521896 271124
rect 521752 235272 521804 235278
rect 521752 235214 521804 235220
rect 521856 231130 521884 271118
rect 521948 247722 521976 276014
rect 522040 271182 522068 346258
rect 523052 326398 523080 436222
rect 523132 417444 523184 417450
rect 523132 417386 523184 417392
rect 523144 351898 523172 417386
rect 523224 414112 523276 414118
rect 523224 414054 523276 414060
rect 523236 380186 523264 414054
rect 523224 380180 523276 380186
rect 523224 380122 523276 380128
rect 523132 351892 523184 351898
rect 523132 351834 523184 351840
rect 523144 350606 523172 351834
rect 523132 350600 523184 350606
rect 523132 350542 523184 350548
rect 523236 346390 523264 380122
rect 523224 346384 523276 346390
rect 523224 346326 523276 346332
rect 523040 326392 523092 326398
rect 523040 326334 523092 326340
rect 522304 302592 522356 302598
rect 522304 302534 522356 302540
rect 522028 271176 522080 271182
rect 522028 271118 522080 271124
rect 521936 247716 521988 247722
rect 521936 247658 521988 247664
rect 521844 231124 521896 231130
rect 521844 231066 521896 231072
rect 521660 224936 521712 224942
rect 521660 224878 521712 224884
rect 521856 219434 521884 231066
rect 521764 219406 521884 219434
rect 521764 202842 521792 219406
rect 521948 216646 521976 247658
rect 522028 235272 522080 235278
rect 522028 235214 522080 235220
rect 522040 219366 522068 235214
rect 522028 219360 522080 219366
rect 522028 219302 522080 219308
rect 521936 216640 521988 216646
rect 521936 216582 521988 216588
rect 521752 202836 521804 202842
rect 521752 202778 521804 202784
rect 522316 193186 522344 302534
rect 523052 293894 523080 326334
rect 524432 295186 524460 437514
rect 525800 436212 525852 436218
rect 525800 436154 525852 436160
rect 524512 433492 524564 433498
rect 524512 433434 524564 433440
rect 524524 315314 524552 433434
rect 524788 425740 524840 425746
rect 524788 425682 524840 425688
rect 524604 414044 524656 414050
rect 524604 413986 524656 413992
rect 524616 347750 524644 413986
rect 524696 413296 524748 413302
rect 524696 413238 524748 413244
rect 524604 347744 524656 347750
rect 524604 347686 524656 347692
rect 524708 343602 524736 413238
rect 524800 369850 524828 425682
rect 524788 369844 524840 369850
rect 524788 369786 524840 369792
rect 524788 350600 524840 350606
rect 524788 350542 524840 350548
rect 524696 343596 524748 343602
rect 524696 343538 524748 343544
rect 524512 315308 524564 315314
rect 524512 315250 524564 315256
rect 524420 295180 524472 295186
rect 524420 295122 524472 295128
rect 523040 293888 523092 293894
rect 523040 293830 523092 293836
rect 524524 289678 524552 315250
rect 524512 289672 524564 289678
rect 524512 289614 524564 289620
rect 524512 281580 524564 281586
rect 524512 281522 524564 281528
rect 523132 278860 523184 278866
rect 523132 278802 523184 278808
rect 523040 270224 523092 270230
rect 523040 270166 523092 270172
rect 523052 200054 523080 270166
rect 523144 238066 523172 278802
rect 524420 278792 524472 278798
rect 524420 278734 524472 278740
rect 523132 238060 523184 238066
rect 523132 238002 523184 238008
rect 523144 220794 523172 238002
rect 524432 222154 524460 278734
rect 524524 226302 524552 281522
rect 524800 273222 524828 350542
rect 525064 302456 525116 302462
rect 525064 302398 525116 302404
rect 524788 273216 524840 273222
rect 524788 273158 524840 273164
rect 524604 271244 524656 271250
rect 524604 271186 524656 271192
rect 524616 228410 524644 271186
rect 524604 228404 524656 228410
rect 524604 228346 524656 228352
rect 524512 226296 524564 226302
rect 524512 226238 524564 226244
rect 524420 222148 524472 222154
rect 524420 222090 524472 222096
rect 523132 220788 523184 220794
rect 523132 220730 523184 220736
rect 524616 204270 524644 228346
rect 524604 204264 524656 204270
rect 524604 204206 524656 204212
rect 523040 200048 523092 200054
rect 523040 199990 523092 199996
rect 522304 193180 522356 193186
rect 522304 193122 522356 193128
rect 520924 153196 520976 153202
rect 520924 153138 520976 153144
rect 518900 153060 518952 153066
rect 518900 153002 518952 153008
rect 518164 139392 518216 139398
rect 518164 139334 518216 139340
rect 517482 124222 517560 124250
rect 517426 124199 517482 124208
rect 516508 124160 516560 124166
rect 516508 124102 516560 124108
rect 514116 123752 514168 123758
rect 514116 123694 514168 123700
rect 514024 122732 514076 122738
rect 514024 122674 514076 122680
rect 508872 122664 508924 122670
rect 508872 122606 508924 122612
rect 502984 99408 503036 99414
rect 502984 99350 503036 99356
rect 423772 99204 423824 99210
rect 423772 99146 423824 99152
rect 374000 98592 374052 98598
rect 374000 98534 374052 98540
rect 345664 98524 345716 98530
rect 345664 98466 345716 98472
rect 336004 98456 336056 98462
rect 336004 98398 336056 98404
rect 322204 97980 322256 97986
rect 322204 97922 322256 97928
rect 320180 94172 320232 94178
rect 320180 94114 320232 94120
rect 317420 90092 317472 90098
rect 317420 90034 317472 90040
rect 316684 73160 316736 73166
rect 316684 73102 316736 73108
rect 316132 72480 316184 72486
rect 316132 72422 316184 72428
rect 316144 16574 316172 72422
rect 316144 16546 316264 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 315028 2984 315080 2990
rect 315028 2926 315080 2932
rect 315040 480 315068 2926
rect 316236 480 316264 16546
rect 317432 6914 317460 90034
rect 318064 85468 318116 85474
rect 318064 85410 318116 85416
rect 318076 16574 318104 85410
rect 320192 16574 320220 94114
rect 318076 16546 318196 16574
rect 320192 16546 320496 16574
rect 317432 6886 318104 6914
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 318076 490 318104 6886
rect 318168 3398 318196 16546
rect 318156 3392 318208 3398
rect 318156 3334 318208 3340
rect 319720 3392 319772 3398
rect 319720 3334 319772 3340
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 3334
rect 320468 490 320496 16546
rect 322112 10668 322164 10674
rect 322112 10610 322164 10616
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 10610
rect 322216 3874 322244 97922
rect 327724 97912 327776 97918
rect 327724 97854 327776 97860
rect 323584 97232 323636 97238
rect 323584 97174 323636 97180
rect 323596 15910 323624 97174
rect 324964 96620 325016 96626
rect 324964 96562 325016 96568
rect 322940 15904 322992 15910
rect 322940 15846 322992 15852
rect 323584 15904 323636 15910
rect 323584 15846 323636 15852
rect 322204 3868 322256 3874
rect 322204 3810 322256 3816
rect 322952 490 322980 15846
rect 324320 10600 324372 10606
rect 324320 10542 324372 10548
rect 324332 3398 324360 10542
rect 324412 6656 324464 6662
rect 324412 6598 324464 6604
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 6598
rect 324976 3330 325004 96562
rect 327736 3738 327764 97854
rect 331220 94376 331272 94382
rect 331220 94318 331272 94324
rect 328460 91656 328512 91662
rect 328460 91598 328512 91604
rect 328472 16574 328500 91598
rect 329840 86216 329892 86222
rect 329840 86158 329892 86164
rect 329852 16574 329880 86158
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 328000 6588 328052 6594
rect 328000 6530 328052 6536
rect 327724 3732 327776 3738
rect 327724 3674 327776 3680
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324964 3324 325016 3330
rect 324964 3266 325016 3272
rect 325620 480 325648 3334
rect 326804 3324 326856 3330
rect 326804 3266 326856 3272
rect 326816 480 326844 3266
rect 328012 480 328040 6530
rect 328748 490 328776 16546
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 331232 490 331260 94318
rect 333980 92948 334032 92954
rect 333980 92890 334032 92896
rect 331864 88868 331916 88874
rect 331864 88810 331916 88816
rect 331876 3398 331904 88810
rect 333992 16574 334020 92890
rect 335360 90160 335412 90166
rect 335360 90102 335412 90108
rect 335372 16574 335400 90102
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 333888 13524 333940 13530
rect 333888 13466 333940 13472
rect 331864 3392 331916 3398
rect 331864 3334 331916 3340
rect 332692 3392 332744 3398
rect 332692 3334 332744 3340
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 3334
rect 333900 480 333928 13466
rect 334636 490 334664 16546
rect 335924 3210 335952 16546
rect 336016 3398 336044 98398
rect 340880 93084 340932 93090
rect 340880 93026 340932 93032
rect 338120 93016 338172 93022
rect 338120 92958 338172 92964
rect 338132 16574 338160 92958
rect 339500 90228 339552 90234
rect 339500 90170 339552 90176
rect 338132 16546 338712 16574
rect 336004 3392 336056 3398
rect 336004 3334 336056 3340
rect 337476 3392 337528 3398
rect 337476 3334 337528 3340
rect 335924 3182 336320 3210
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3182
rect 337488 480 337516 3334
rect 338684 480 338712 16546
rect 339512 490 339540 90170
rect 340892 3398 340920 93026
rect 342260 88936 342312 88942
rect 342260 88878 342312 88884
rect 340972 85400 341024 85406
rect 340972 85342 341024 85348
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 85342
rect 342272 6914 342300 88878
rect 342904 85332 342956 85338
rect 342904 85274 342956 85280
rect 342916 16574 342944 85274
rect 342916 16546 343036 16574
rect 342272 6886 342944 6914
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 342916 490 342944 6886
rect 343008 3398 343036 16546
rect 345676 3398 345704 98466
rect 352564 97844 352616 97850
rect 352564 97786 352616 97792
rect 346400 89684 346452 89690
rect 346400 89626 346452 89632
rect 346412 16574 346440 89626
rect 346412 16546 346992 16574
rect 345756 6520 345808 6526
rect 345756 6462 345808 6468
rect 342996 3392 343048 3398
rect 342996 3334 343048 3340
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 345664 3392 345716 3398
rect 345664 3334 345716 3340
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3334
rect 345768 480 345796 6462
rect 346964 480 346992 16546
rect 352576 6458 352604 97786
rect 359464 97776 359516 97782
rect 359464 97718 359516 97724
rect 353944 94444 353996 94450
rect 353944 94386 353996 94392
rect 353300 91724 353352 91730
rect 353300 91666 353352 91672
rect 353312 16574 353340 91666
rect 353312 16546 353616 16574
rect 352840 6588 352892 6594
rect 352840 6530 352892 6536
rect 352564 6452 352616 6458
rect 352564 6394 352616 6400
rect 351644 3936 351696 3942
rect 351644 3878 351696 3884
rect 349252 3800 349304 3806
rect 349252 3742 349304 3748
rect 348056 3392 348108 3398
rect 348056 3334 348108 3340
rect 348068 480 348096 3334
rect 349264 480 349292 3742
rect 350448 3664 350500 3670
rect 350448 3606 350500 3612
rect 350460 480 350488 3606
rect 351656 480 351684 3878
rect 352852 480 352880 6530
rect 353588 490 353616 16546
rect 353956 4146 353984 94386
rect 356704 90296 356756 90302
rect 356704 90238 356756 90244
rect 356336 6520 356388 6526
rect 356336 6462 356388 6468
rect 353944 4140 353996 4146
rect 353944 4082 353996 4088
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 353864 598 354076 626
rect 353864 490 353892 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 462 353892 490
rect 354048 480 354076 598
rect 355244 480 355272 4082
rect 356348 480 356376 6462
rect 356716 3670 356744 90238
rect 357440 87576 357492 87582
rect 357440 87518 357492 87524
rect 357452 6914 357480 87518
rect 357532 83904 357584 83910
rect 357532 83846 357584 83852
rect 357544 11694 357572 83846
rect 357532 11688 357584 11694
rect 357532 11630 357584 11636
rect 358728 11688 358780 11694
rect 358728 11630 358780 11636
rect 357452 6886 357572 6914
rect 356704 3664 356756 3670
rect 356704 3606 356756 3612
rect 357544 480 357572 6886
rect 358740 480 358768 11630
rect 359476 6322 359504 97718
rect 363604 97708 363656 97714
rect 363604 97650 363656 97656
rect 360844 93832 360896 93838
rect 360844 93774 360896 93780
rect 360200 88324 360252 88330
rect 360200 88266 360252 88272
rect 360212 16574 360240 88266
rect 360212 16546 360792 16574
rect 359924 6384 359976 6390
rect 359924 6326 359976 6332
rect 359464 6316 359516 6322
rect 359464 6258 359516 6264
rect 359936 480 359964 6326
rect 360764 3210 360792 16546
rect 360856 3398 360884 93774
rect 362316 9104 362368 9110
rect 362316 9046 362368 9052
rect 360844 3392 360896 3398
rect 360844 3334 360896 3340
rect 360764 3182 361160 3210
rect 361132 480 361160 3182
rect 362328 480 362356 9046
rect 363616 5166 363644 97650
rect 370504 97640 370556 97646
rect 370504 97582 370556 97588
rect 369124 97572 369176 97578
rect 369124 97514 369176 97520
rect 364984 93764 365036 93770
rect 364984 93706 365036 93712
rect 364340 88256 364392 88262
rect 364340 88198 364392 88204
rect 364352 16574 364380 88198
rect 364352 16546 364656 16574
rect 363604 5160 363656 5166
rect 363604 5102 363656 5108
rect 363512 3392 363564 3398
rect 363512 3334 363564 3340
rect 363524 480 363552 3334
rect 364628 480 364656 16546
rect 364996 3058 365024 93706
rect 367744 93696 367796 93702
rect 367744 93638 367796 93644
rect 367100 86896 367152 86902
rect 367100 86838 367152 86844
rect 365812 83836 365864 83842
rect 365812 83778 365864 83784
rect 364984 3052 365036 3058
rect 364984 2994 365036 3000
rect 365824 480 365852 83778
rect 367112 6914 367140 86838
rect 367756 16574 367784 93638
rect 367756 16546 367876 16574
rect 367112 6886 367784 6914
rect 367008 3052 367060 3058
rect 367008 2994 367060 3000
rect 367020 480 367048 2994
rect 367756 490 367784 6886
rect 367848 3398 367876 16546
rect 367836 3392 367888 3398
rect 367836 3334 367888 3340
rect 369136 3058 369164 97514
rect 370516 5234 370544 97582
rect 374012 6914 374040 98534
rect 413284 98388 413336 98394
rect 413284 98330 413336 98336
rect 374644 93628 374696 93634
rect 374644 93570 374696 93576
rect 374092 88188 374144 88194
rect 374092 88130 374144 88136
rect 374104 16574 374132 88130
rect 374104 16546 374592 16574
rect 374012 6886 374132 6914
rect 370504 5228 370556 5234
rect 370504 5170 370556 5176
rect 372896 5092 372948 5098
rect 372896 5034 372948 5040
rect 369400 3664 369452 3670
rect 369400 3606 369452 3612
rect 369124 3052 369176 3058
rect 369124 2994 369176 3000
rect 368032 598 368244 626
rect 368032 490 368060 598
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 462 368060 490
rect 368216 480 368244 598
rect 369412 480 369440 3606
rect 370596 3392 370648 3398
rect 370596 3334 370648 3340
rect 370608 480 370636 3334
rect 371700 3052 371752 3058
rect 371700 2994 371752 3000
rect 371712 480 371740 2994
rect 372908 480 372936 5034
rect 374104 480 374132 6886
rect 374564 3210 374592 16546
rect 374656 3398 374684 93570
rect 378784 92472 378836 92478
rect 378784 92414 378836 92420
rect 378140 88120 378192 88126
rect 378140 88062 378192 88068
rect 375380 85264 375432 85270
rect 375380 85206 375432 85212
rect 375392 16574 375420 85206
rect 377404 82408 377456 82414
rect 377404 82350 377456 82356
rect 375392 16546 376064 16574
rect 374644 3392 374696 3398
rect 374644 3334 374696 3340
rect 374564 3182 375328 3210
rect 375300 480 375328 3182
rect 376036 490 376064 16546
rect 377416 3058 377444 82350
rect 378152 16574 378180 88062
rect 378152 16546 378456 16574
rect 377680 3392 377732 3398
rect 377680 3334 377732 3340
rect 377404 3052 377456 3058
rect 377404 2994 377456 3000
rect 376312 598 376524 626
rect 376312 490 376340 598
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 462 376340 490
rect 376496 480 376524 598
rect 377692 480 377720 3334
rect 378428 490 378456 16546
rect 378796 3398 378824 92414
rect 382924 92404 382976 92410
rect 382924 92346 382976 92352
rect 381544 86828 381596 86834
rect 381544 86770 381596 86776
rect 381556 3806 381584 86770
rect 382372 86760 382424 86766
rect 382372 86702 382424 86708
rect 381544 3800 381596 3806
rect 381544 3742 381596 3748
rect 378784 3392 378836 3398
rect 378784 3334 378836 3340
rect 381176 3392 381228 3398
rect 381176 3334 381228 3340
rect 379980 3052 380032 3058
rect 379980 2994 380032 3000
rect 378704 598 378916 626
rect 378704 490 378732 598
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 462 378732 490
rect 378888 480 378916 598
rect 379992 480 380020 2994
rect 381188 480 381216 3334
rect 382384 480 382412 86702
rect 382936 3398 382964 92346
rect 387800 92336 387852 92342
rect 387800 92278 387852 92284
rect 385684 89616 385736 89622
rect 385684 89558 385736 89564
rect 385592 12300 385644 12306
rect 385592 12242 385644 12248
rect 383568 3868 383620 3874
rect 383568 3810 383620 3816
rect 382924 3392 382976 3398
rect 382924 3334 382976 3340
rect 383580 480 383608 3810
rect 384764 3392 384816 3398
rect 384764 3334 384816 3340
rect 384776 480 384804 3334
rect 385604 3074 385632 12242
rect 385696 3262 385724 89558
rect 385684 3256 385736 3262
rect 385684 3198 385736 3204
rect 387156 3256 387208 3262
rect 387156 3198 387208 3204
rect 385604 3046 386000 3074
rect 385972 480 386000 3046
rect 387168 480 387196 3198
rect 387812 490 387840 92278
rect 389824 92268 389876 92274
rect 389824 92210 389876 92216
rect 389456 12232 389508 12238
rect 389456 12174 389508 12180
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 12174
rect 389836 3398 389864 92210
rect 407764 91044 407816 91050
rect 407764 90986 407816 90992
rect 403624 90976 403676 90982
rect 403624 90918 403676 90924
rect 392584 88052 392636 88058
rect 392584 87994 392636 88000
rect 392596 16574 392624 87994
rect 395344 86692 395396 86698
rect 395344 86634 395396 86640
rect 393964 82272 394016 82278
rect 393964 82214 394016 82220
rect 392596 16546 392716 16574
rect 392584 12164 392636 12170
rect 392584 12106 392636 12112
rect 390652 3732 390704 3738
rect 390652 3674 390704 3680
rect 389824 3392 389876 3398
rect 389824 3334 389876 3340
rect 390664 480 390692 3674
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 392596 490 392624 12106
rect 392688 4010 392716 16546
rect 392676 4004 392728 4010
rect 392676 3946 392728 3952
rect 393976 3874 394004 82214
rect 395252 8084 395304 8090
rect 395252 8026 395304 8032
rect 394240 4004 394292 4010
rect 394240 3946 394292 3952
rect 393964 3868 394016 3874
rect 393964 3810 394016 3816
rect 392872 598 393084 626
rect 392872 490 392900 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 462 392900 490
rect 393056 480 393084 598
rect 394252 480 394280 3946
rect 395264 3482 395292 8026
rect 395356 3670 395384 86634
rect 400220 82476 400272 82482
rect 400220 82418 400272 82424
rect 396724 82340 396776 82346
rect 396724 82282 396776 82288
rect 396080 12096 396132 12102
rect 396080 12038 396132 12044
rect 395344 3664 395396 3670
rect 395344 3606 395396 3612
rect 395264 3454 395384 3482
rect 395356 480 395384 3454
rect 396092 490 396120 12038
rect 396736 3738 396764 82282
rect 399484 80844 399536 80850
rect 399484 80786 399536 80792
rect 398840 12028 398892 12034
rect 398840 11970 398892 11976
rect 396724 3732 396776 3738
rect 396724 3674 396776 3680
rect 397736 3664 397788 3670
rect 397736 3606 397788 3612
rect 396368 598 396580 626
rect 396368 490 396396 598
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 462 396396 490
rect 396552 480 396580 598
rect 397748 480 397776 3606
rect 398852 3398 398880 11970
rect 398932 8016 398984 8022
rect 398932 7958 398984 7964
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 7958
rect 399496 3670 399524 80786
rect 400232 16574 400260 82418
rect 400232 16546 400904 16574
rect 399484 3664 399536 3670
rect 399484 3606 399536 3612
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 400876 490 400904 16546
rect 403532 11960 403584 11966
rect 403532 11902 403584 11908
rect 402520 7948 402572 7954
rect 402520 7890 402572 7896
rect 401152 598 401364 626
rect 401152 490 401180 598
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 462 401180 490
rect 401336 480 401364 598
rect 402532 480 402560 7890
rect 403544 3210 403572 11902
rect 403636 3398 403664 90918
rect 406384 86624 406436 86630
rect 406384 86566 406436 86572
rect 404360 15904 404412 15910
rect 404360 15846 404412 15852
rect 403624 3392 403676 3398
rect 403624 3334 403676 3340
rect 403544 3182 403664 3210
rect 403636 480 403664 3182
rect 404372 490 404400 15846
rect 406016 7880 406068 7886
rect 406016 7822 406068 7828
rect 404648 598 404860 626
rect 404648 490 404676 598
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 462 404676 490
rect 404832 480 404860 598
rect 406028 480 406056 7822
rect 406396 4078 406424 86566
rect 407212 11892 407264 11898
rect 407212 11834 407264 11840
rect 406384 4072 406436 4078
rect 406384 4014 406436 4020
rect 407224 480 407252 11834
rect 407776 3942 407804 90986
rect 410524 89548 410576 89554
rect 410524 89490 410576 89496
rect 410432 11824 410484 11830
rect 410432 11766 410484 11772
rect 409604 7812 409656 7818
rect 409604 7754 409656 7760
rect 407764 3936 407816 3942
rect 407764 3878 407816 3884
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 409616 480 409644 7754
rect 410444 3482 410472 11766
rect 410536 4146 410564 89490
rect 411904 80776 411956 80782
rect 411904 80718 411956 80724
rect 411916 16574 411944 80718
rect 411916 16546 412036 16574
rect 410524 4140 410576 4146
rect 410524 4082 410576 4088
rect 412008 3806 412036 16546
rect 413100 7744 413152 7750
rect 413100 7686 413152 7692
rect 411904 3800 411956 3806
rect 411904 3742 411956 3748
rect 411996 3800 412048 3806
rect 411996 3742 412048 3748
rect 410444 3454 410840 3482
rect 410812 480 410840 3454
rect 411916 480 411944 3742
rect 413112 480 413140 7686
rect 413296 3126 413324 98330
rect 414664 98320 414716 98326
rect 414664 98262 414716 98268
rect 414296 11756 414348 11762
rect 414296 11698 414348 11704
rect 413284 3120 413336 3126
rect 413284 3062 413336 3068
rect 414308 480 414336 11698
rect 414676 3398 414704 98262
rect 416780 93560 416832 93566
rect 416780 93502 416832 93508
rect 416792 16574 416820 93502
rect 421564 93492 421616 93498
rect 421564 93434 421616 93440
rect 418804 83768 418856 83774
rect 418804 83710 418856 83716
rect 416792 16546 417464 16574
rect 416688 7676 416740 7682
rect 416688 7618 416740 7624
rect 415492 5024 415544 5030
rect 415492 4966 415544 4972
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 4966
rect 416700 480 416728 7618
rect 417436 490 417464 16546
rect 418816 4078 418844 83710
rect 418988 6452 419040 6458
rect 418988 6394 419040 6400
rect 418804 4072 418856 4078
rect 418804 4014 418856 4020
rect 417712 598 417924 626
rect 417712 490 417740 598
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 462 417740 490
rect 417896 480 417924 598
rect 419000 480 419028 6394
rect 421576 3398 421604 93434
rect 422576 3868 422628 3874
rect 422576 3810 422628 3816
rect 421380 3392 421432 3398
rect 421380 3334 421432 3340
rect 421564 3392 421616 3398
rect 421564 3334 421616 3340
rect 420184 3120 420236 3126
rect 420184 3062 420236 3068
rect 420196 480 420224 3062
rect 421392 480 421420 3334
rect 422588 480 422616 3810
rect 423784 480 423812 99146
rect 435364 99136 435416 99142
rect 435364 99078 435416 99084
rect 425704 97504 425756 97510
rect 425704 97446 425756 97452
rect 425716 6322 425744 97446
rect 429844 97436 429896 97442
rect 429844 97378 429896 97384
rect 427820 87984 427872 87990
rect 427820 87926 427872 87932
rect 427832 16574 427860 87926
rect 427832 16546 428504 16574
rect 426164 6384 426216 6390
rect 426164 6326 426216 6332
rect 425704 6316 425756 6322
rect 425704 6258 425756 6264
rect 424968 4140 425020 4146
rect 424968 4082 425020 4088
rect 424980 480 425008 4082
rect 426176 480 426204 6326
rect 427268 3392 427320 3398
rect 427268 3334 427320 3340
rect 427280 480 427308 3334
rect 428476 480 428504 16546
rect 429660 5160 429712 5166
rect 429660 5102 429712 5108
rect 429672 480 429700 5102
rect 429856 5098 429884 97378
rect 430580 92200 430632 92206
rect 430580 92142 430632 92148
rect 430592 16574 430620 92142
rect 432604 92132 432656 92138
rect 432604 92074 432656 92080
rect 430592 16546 430896 16574
rect 429844 5092 429896 5098
rect 429844 5034 429896 5040
rect 430868 480 430896 16546
rect 432052 4004 432104 4010
rect 432052 3946 432104 3952
rect 432064 480 432092 3946
rect 432616 3398 432644 92074
rect 433248 5228 433300 5234
rect 433248 5170 433300 5176
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 433260 480 433288 5170
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 434456 480 434484 3334
rect 435376 3058 435404 99078
rect 440884 99068 440936 99074
rect 440884 99010 440936 99016
rect 436744 97368 436796 97374
rect 436744 97310 436796 97316
rect 436756 16574 436784 97310
rect 438860 87916 438912 87922
rect 438860 87858 438912 87864
rect 438872 16574 438900 87858
rect 436756 16546 436876 16574
rect 438872 16546 439176 16574
rect 436744 4072 436796 4078
rect 436744 4014 436796 4020
rect 435548 3936 435600 3942
rect 435548 3878 435600 3884
rect 435364 3052 435416 3058
rect 435364 2994 435416 3000
rect 435560 480 435588 3878
rect 436756 480 436784 4014
rect 436848 4010 436876 16546
rect 436836 4004 436888 4010
rect 436836 3946 436888 3952
rect 437940 3052 437992 3058
rect 437940 2994 437992 3000
rect 437952 480 437980 2994
rect 439148 480 439176 16546
rect 440896 3874 440924 99010
rect 457444 99000 457496 99006
rect 457444 98942 457496 98948
rect 450542 97472 450598 97481
rect 450542 97407 450598 97416
rect 447782 97336 447838 97345
rect 443644 97300 443696 97306
rect 447782 97271 447838 97280
rect 443644 97242 443696 97248
rect 442264 89480 442316 89486
rect 442264 89422 442316 89428
rect 441620 86556 441672 86562
rect 441620 86498 441672 86504
rect 441632 16574 441660 86498
rect 441632 16546 442212 16574
rect 441528 7608 441580 7614
rect 441528 7550 441580 7556
rect 440884 3868 440936 3874
rect 440884 3810 440936 3816
rect 440332 3800 440384 3806
rect 440332 3742 440384 3748
rect 440344 480 440372 3742
rect 441540 480 441568 7550
rect 442184 3210 442212 16546
rect 442276 3398 442304 89422
rect 443656 3806 443684 97242
rect 446404 92064 446456 92070
rect 446404 92006 446456 92012
rect 445024 3868 445076 3874
rect 445024 3810 445076 3816
rect 443644 3800 443696 3806
rect 443644 3742 443696 3748
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 442264 3392 442316 3398
rect 442264 3334 442316 3340
rect 442184 3182 442672 3210
rect 442644 480 442672 3182
rect 443840 480 443868 3674
rect 445036 480 445064 3810
rect 446220 3392 446272 3398
rect 446220 3334 446272 3340
rect 446232 480 446260 3334
rect 446416 2990 446444 92006
rect 447796 6322 447824 97271
rect 448520 93424 448572 93430
rect 448520 93366 448572 93372
rect 447416 6316 447468 6322
rect 447416 6258 447468 6264
rect 447784 6316 447836 6322
rect 447784 6258 447836 6264
rect 446404 2984 446456 2990
rect 446404 2926 446456 2932
rect 447428 480 447456 6258
rect 448532 2774 448560 93366
rect 448612 86488 448664 86494
rect 448612 86430 448664 86436
rect 448624 7614 448652 86430
rect 448612 7608 448664 7614
rect 448612 7550 448664 7556
rect 449808 7608 449860 7614
rect 449808 7550 449860 7556
rect 449164 3528 449216 3534
rect 449164 3470 449216 3476
rect 449176 3398 449204 3470
rect 449164 3392 449216 3398
rect 449164 3334 449216 3340
rect 448532 2746 448652 2774
rect 448624 480 448652 2746
rect 449820 480 449848 7550
rect 450556 5030 450584 97407
rect 454684 95192 454736 95198
rect 454684 95134 454736 95140
rect 453304 91996 453356 92002
rect 453304 91938 453356 91944
rect 453212 13456 453264 13462
rect 453212 13398 453264 13404
rect 450544 5024 450596 5030
rect 450544 4966 450596 4972
rect 450912 3664 450964 3670
rect 450912 3606 450964 3612
rect 450924 480 450952 3606
rect 452108 2984 452160 2990
rect 452108 2926 452160 2932
rect 452120 480 452148 2926
rect 453224 2774 453252 13398
rect 453316 4146 453344 91938
rect 454500 5092 454552 5098
rect 454500 5034 454552 5040
rect 453304 4140 453356 4146
rect 453304 4082 453356 4088
rect 453224 2746 453344 2774
rect 453316 480 453344 2746
rect 454512 480 454540 5034
rect 454696 3670 454724 95134
rect 456892 13388 456944 13394
rect 456892 13330 456944 13336
rect 455696 4140 455748 4146
rect 455696 4082 455748 4088
rect 454684 3664 454736 3670
rect 454684 3606 454736 3612
rect 455708 480 455736 4082
rect 456904 480 456932 13330
rect 457456 3534 457484 98942
rect 458180 98932 458232 98938
rect 458180 98874 458232 98880
rect 458192 16574 458220 98874
rect 467104 98864 467156 98870
rect 467104 98806 467156 98812
rect 461584 96552 461636 96558
rect 461584 96494 461636 96500
rect 460204 91928 460256 91934
rect 460204 91870 460256 91876
rect 458192 16546 459232 16574
rect 457444 3528 457496 3534
rect 457444 3470 457496 3476
rect 458088 3256 458140 3262
rect 458088 3198 458140 3204
rect 458100 480 458128 3198
rect 459204 480 459232 16546
rect 459928 13320 459980 13326
rect 459928 13262 459980 13268
rect 459940 490 459968 13262
rect 460216 4146 460244 91870
rect 461596 16574 461624 96494
rect 464344 95124 464396 95130
rect 464344 95066 464396 95072
rect 461596 16546 461716 16574
rect 460204 4140 460256 4146
rect 460204 4082 460256 4088
rect 461584 3868 461636 3874
rect 461584 3810 461636 3816
rect 460216 598 460428 626
rect 460216 490 460244 598
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 462 460244 490
rect 460400 480 460428 598
rect 461596 480 461624 3810
rect 461688 3806 461716 16546
rect 463976 13252 464028 13258
rect 463976 13194 464028 13200
rect 462780 4140 462832 4146
rect 462780 4082 462832 4088
rect 461676 3800 461728 3806
rect 461676 3742 461728 3748
rect 462792 480 462820 4082
rect 463988 480 464016 13194
rect 464356 4078 464384 95066
rect 465724 91860 465776 91866
rect 465724 91802 465776 91808
rect 465172 90840 465224 90846
rect 465172 90782 465224 90788
rect 465184 16574 465212 90782
rect 465184 16546 465672 16574
rect 464344 4072 464396 4078
rect 464344 4014 464396 4020
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 465184 480 465212 3538
rect 465644 626 465672 16546
rect 465736 3330 465764 91802
rect 467116 3602 467144 98806
rect 490564 98796 490616 98802
rect 490564 98738 490616 98744
rect 468484 96484 468536 96490
rect 468484 96426 468536 96432
rect 468496 3874 468524 96426
rect 472624 96416 472676 96422
rect 472624 96358 472676 96364
rect 471244 90908 471296 90914
rect 471244 90850 471296 90856
rect 470600 86420 470652 86426
rect 470600 86362 470652 86368
rect 468484 3868 468536 3874
rect 468484 3810 468536 3816
rect 468668 3732 468720 3738
rect 468668 3674 468720 3680
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 465724 3324 465776 3330
rect 465724 3266 465776 3272
rect 467472 3324 467524 3330
rect 467472 3266 467524 3272
rect 465644 598 465856 626
rect 465828 490 465856 598
rect 466104 598 466316 626
rect 466104 490 466132 598
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 462 466132 490
rect 466288 480 466316 598
rect 467484 480 467512 3266
rect 468680 480 468708 3674
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 470612 490 470640 86362
rect 471256 3602 471284 90850
rect 472256 6248 472308 6254
rect 472256 6190 472308 6196
rect 471244 3596 471296 3602
rect 471244 3538 471296 3544
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 6190
rect 472636 3942 472664 96358
rect 475384 96348 475436 96354
rect 475384 96290 475436 96296
rect 472716 85196 472768 85202
rect 472716 85138 472768 85144
rect 472624 3936 472676 3942
rect 472624 3878 472676 3884
rect 472728 2922 472756 85138
rect 473452 4072 473504 4078
rect 473452 4014 473504 4020
rect 472716 2916 472768 2922
rect 472716 2858 472768 2864
rect 473464 480 473492 4014
rect 475396 3738 475424 96290
rect 479524 96280 479576 96286
rect 479524 96222 479576 96228
rect 476764 90772 476816 90778
rect 476764 90714 476816 90720
rect 475752 6316 475804 6322
rect 475752 6258 475804 6264
rect 475384 3732 475436 3738
rect 475384 3674 475436 3680
rect 474556 2916 474608 2922
rect 474556 2858 474608 2864
rect 474568 480 474596 2858
rect 475764 480 475792 6258
rect 476776 4010 476804 90714
rect 478144 13184 478196 13190
rect 478144 13126 478196 13132
rect 476948 9036 477000 9042
rect 476948 8978 477000 8984
rect 476764 4004 476816 4010
rect 476764 3946 476816 3952
rect 476960 480 476988 8978
rect 478156 480 478184 13126
rect 479536 4146 479564 96222
rect 483020 96212 483072 96218
rect 483020 96154 483072 96160
rect 482284 85128 482336 85134
rect 482284 85070 482336 85076
rect 482192 13116 482244 13122
rect 482192 13058 482244 13064
rect 481732 8968 481784 8974
rect 481732 8910 481784 8916
rect 479524 4140 479576 4146
rect 479524 4082 479576 4088
rect 480536 4140 480588 4146
rect 480536 4082 480588 4088
rect 479340 3460 479392 3466
rect 479340 3402 479392 3408
rect 479352 480 479380 3402
rect 480548 480 480576 4082
rect 481744 480 481772 8910
rect 482204 626 482232 13058
rect 482296 3330 482324 85070
rect 483032 16574 483060 96154
rect 485044 95056 485096 95062
rect 485044 94998 485096 95004
rect 483032 16546 484072 16574
rect 482284 3324 482336 3330
rect 482284 3266 482336 3272
rect 482204 598 482416 626
rect 482388 490 482416 598
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 16546
rect 485056 3398 485084 94998
rect 489184 94988 489236 94994
rect 489184 94930 489236 94936
rect 486424 90704 486476 90710
rect 486424 90646 486476 90652
rect 485228 4004 485280 4010
rect 485228 3946 485280 3952
rect 485044 3392 485096 3398
rect 485044 3334 485096 3340
rect 485240 480 485268 3946
rect 486436 3466 486464 90646
rect 489196 3738 489224 94930
rect 490012 19984 490064 19990
rect 490012 19926 490064 19932
rect 490024 6914 490052 19926
rect 489932 6886 490052 6914
rect 487620 3732 487672 3738
rect 487620 3674 487672 3680
rect 489184 3732 489236 3738
rect 489184 3674 489236 3680
rect 486424 3460 486476 3466
rect 486424 3402 486476 3408
rect 486424 3324 486476 3330
rect 486424 3266 486476 3272
rect 486436 480 486464 3266
rect 487632 480 487660 3674
rect 488816 3460 488868 3466
rect 488816 3402 488868 3408
rect 488828 480 488856 3402
rect 489932 480 489960 6886
rect 490576 3398 490604 98738
rect 494060 96144 494112 96150
rect 494060 96086 494112 96092
rect 493324 90636 493376 90642
rect 493324 90578 493376 90584
rect 492680 85060 492732 85066
rect 492680 85002 492732 85008
rect 492692 16574 492720 85002
rect 492692 16546 493088 16574
rect 491116 3936 491168 3942
rect 491116 3878 491168 3884
rect 490564 3392 490616 3398
rect 490564 3334 490616 3340
rect 491128 480 491156 3878
rect 492312 3392 492364 3398
rect 492312 3334 492364 3340
rect 492324 480 492352 3334
rect 493060 490 493088 16546
rect 493336 2990 493364 90578
rect 494072 16574 494100 96086
rect 500960 96076 501012 96082
rect 500960 96018 501012 96024
rect 497464 90568 497516 90574
rect 497464 90510 497516 90516
rect 496820 86352 496872 86358
rect 496820 86294 496872 86300
rect 496832 16574 496860 86294
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 493324 2984 493376 2990
rect 493324 2926 493376 2932
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 16546
rect 495900 2984 495952 2990
rect 495900 2926 495952 2932
rect 495912 480 495940 2926
rect 497108 480 497136 16546
rect 497476 3398 497504 90510
rect 500224 90500 500276 90506
rect 500224 90442 500276 90448
rect 499580 84992 499632 84998
rect 499580 84934 499632 84940
rect 499592 6914 499620 84934
rect 500236 16574 500264 90442
rect 500972 16574 501000 96018
rect 507860 96008 507912 96014
rect 507860 95950 507912 95956
rect 502984 94920 503036 94926
rect 502984 94862 503036 94868
rect 502996 16574 503024 94862
rect 504364 90432 504416 90438
rect 504364 90374 504416 90380
rect 500236 16546 500356 16574
rect 500972 16546 501368 16574
rect 502996 16546 503116 16574
rect 499592 6886 500264 6914
rect 498200 3868 498252 3874
rect 498200 3810 498252 3816
rect 497464 3392 497516 3398
rect 497464 3334 497516 3340
rect 498212 480 498240 3810
rect 499396 3392 499448 3398
rect 499396 3334 499448 3340
rect 499408 480 499436 3334
rect 500236 3210 500264 6886
rect 500328 3330 500356 16546
rect 500316 3324 500368 3330
rect 500316 3266 500368 3272
rect 500236 3182 500632 3210
rect 500604 480 500632 3182
rect 501340 490 501368 16546
rect 503088 3874 503116 16546
rect 504180 4956 504232 4962
rect 504180 4898 504232 4904
rect 503076 3868 503128 3874
rect 503076 3810 503128 3816
rect 502984 3324 503036 3330
rect 502984 3266 503036 3272
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 3266
rect 504192 480 504220 4898
rect 504376 3058 504404 90374
rect 506480 89412 506532 89418
rect 506480 89354 506532 89360
rect 505376 3800 505428 3806
rect 505376 3742 505428 3748
rect 504364 3052 504416 3058
rect 504364 2994 504416 3000
rect 505388 480 505416 3742
rect 506492 480 506520 89354
rect 506572 24132 506624 24138
rect 506572 24074 506624 24080
rect 506584 16574 506612 24074
rect 507872 16574 507900 95950
rect 518900 95940 518952 95946
rect 518900 95882 518952 95888
rect 512000 94852 512052 94858
rect 512000 94794 512052 94800
rect 511264 89344 511316 89350
rect 511264 89286 511316 89292
rect 510620 83700 510672 83706
rect 510620 83642 510672 83648
rect 510632 16574 510660 83642
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511212 16574
rect 507228 490 507256 16546
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 16546
rect 510068 3052 510120 3058
rect 510068 2994 510120 3000
rect 510080 480 510108 2994
rect 511184 2938 511212 16546
rect 511276 3058 511304 89286
rect 511264 3052 511316 3058
rect 511264 2994 511316 3000
rect 511184 2910 511304 2938
rect 511276 480 511304 2910
rect 512012 490 512040 94794
rect 515404 91792 515456 91798
rect 515404 91734 515456 91740
rect 514852 26920 514904 26926
rect 514852 26862 514904 26868
rect 514864 6914 514892 26862
rect 514772 6886 514892 6914
rect 513564 3052 513616 3058
rect 513564 2994 513616 3000
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 2994
rect 514772 480 514800 6886
rect 515416 3398 515444 91734
rect 518164 89276 518216 89282
rect 518164 89218 518216 89224
rect 517520 83632 517572 83638
rect 517520 83574 517572 83580
rect 517532 16574 517560 83574
rect 517532 16546 517928 16574
rect 515956 3664 516008 3670
rect 515956 3606 516008 3612
rect 515404 3392 515456 3398
rect 515404 3334 515456 3340
rect 515968 480 515996 3606
rect 517152 3392 517204 3398
rect 517152 3334 517204 3340
rect 517164 480 517192 3334
rect 517900 490 517928 16546
rect 518176 4146 518204 89218
rect 518912 16574 518940 95882
rect 520924 94784 520976 94790
rect 520924 94726 520976 94732
rect 518912 16546 519584 16574
rect 518164 4140 518216 4146
rect 518164 4082 518216 4088
rect 518176 598 518388 626
rect 518176 490 518204 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 462 518204 490
rect 518360 480 518388 598
rect 519556 480 519584 16546
rect 520740 4140 520792 4146
rect 520740 4082 520792 4088
rect 520752 480 520780 4082
rect 520936 3602 520964 94726
rect 522304 89208 522356 89214
rect 522304 89150 522356 89156
rect 521660 18624 521712 18630
rect 521660 18566 521712 18572
rect 521672 16574 521700 18566
rect 521672 16546 521884 16574
rect 520924 3596 520976 3602
rect 520924 3538 520976 3544
rect 521856 480 521884 16546
rect 522316 2990 522344 89150
rect 524420 84924 524472 84930
rect 524420 84866 524472 84872
rect 524432 16574 524460 84866
rect 525076 20670 525104 302398
rect 525812 293962 525840 436154
rect 525892 432064 525944 432070
rect 525892 432006 525944 432012
rect 525904 322250 525932 432006
rect 525984 415472 526036 415478
rect 525984 415414 526036 415420
rect 525996 349858 526024 415414
rect 525984 349852 526036 349858
rect 525984 349794 526036 349800
rect 525892 322244 525944 322250
rect 525892 322186 525944 322192
rect 525800 293956 525852 293962
rect 525800 293898 525852 293904
rect 525904 289746 525932 322186
rect 526456 307086 526484 699654
rect 529940 438932 529992 438938
rect 529940 438874 529992 438880
rect 528744 437504 528796 437510
rect 528744 437446 528796 437452
rect 527180 436144 527232 436150
rect 527180 436086 527232 436092
rect 527192 309806 527220 436086
rect 528652 433424 528704 433430
rect 528652 433366 528704 433372
rect 528560 431996 528612 432002
rect 528560 431938 528612 431944
rect 527180 309800 527232 309806
rect 527180 309742 527232 309748
rect 526444 307080 526496 307086
rect 526444 307022 526496 307028
rect 526444 299600 526496 299606
rect 526444 299542 526496 299548
rect 525892 289740 525944 289746
rect 525892 289682 525944 289688
rect 525892 271924 525944 271930
rect 525892 271866 525944 271872
rect 525800 269136 525852 269142
rect 525800 269078 525852 269084
rect 525812 200122 525840 269078
rect 525904 204950 525932 271866
rect 525892 204944 525944 204950
rect 525892 204886 525944 204892
rect 525800 200116 525852 200122
rect 525800 200058 525852 200064
rect 526456 126954 526484 299542
rect 527192 292466 527220 309742
rect 527180 292460 527232 292466
rect 527180 292402 527232 292408
rect 528572 289814 528600 431938
rect 528664 291106 528692 433366
rect 528756 295254 528784 437446
rect 528836 295996 528888 296002
rect 528836 295938 528888 295944
rect 528744 295248 528796 295254
rect 528744 295190 528796 295196
rect 528652 291100 528704 291106
rect 528652 291042 528704 291048
rect 528560 289808 528612 289814
rect 528560 289750 528612 289756
rect 528652 273216 528704 273222
rect 528652 273158 528704 273164
rect 528664 233918 528692 273158
rect 528652 233912 528704 233918
rect 528652 233854 528704 233860
rect 528664 206922 528692 233854
rect 528652 206916 528704 206922
rect 528652 206858 528704 206864
rect 528848 153134 528876 295938
rect 529952 295322 529980 438874
rect 530032 434784 530084 434790
rect 530032 434726 530084 434732
rect 529940 295316 529992 295322
rect 529940 295258 529992 295264
rect 530044 292534 530072 434726
rect 530124 433356 530176 433362
rect 530124 433298 530176 433304
rect 530032 292528 530084 292534
rect 530032 292470 530084 292476
rect 530136 291174 530164 433298
rect 558932 304706 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 324358 579660 325207
rect 579620 324352 579672 324358
rect 579620 324294 579672 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 558920 304700 558972 304706
rect 558920 304642 558972 304648
rect 580276 304638 580304 577623
rect 580354 564360 580410 564369
rect 580354 564295 580410 564304
rect 580264 304632 580316 304638
rect 580264 304574 580316 304580
rect 580368 304570 580396 564295
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580356 304564 580408 304570
rect 580356 304506 580408 304512
rect 580460 304434 580488 431559
rect 580538 418296 580594 418305
rect 580538 418231 580594 418240
rect 580552 304502 580580 418231
rect 580630 365120 580686 365129
rect 580630 365055 580686 365064
rect 580540 304496 580592 304502
rect 580540 304438 580592 304444
rect 580448 304428 580500 304434
rect 580448 304370 580500 304376
rect 580644 304366 580672 365055
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580632 304360 580684 304366
rect 580632 304302 580684 304308
rect 580736 304298 580764 351863
rect 582392 305726 582420 511255
rect 582470 484664 582526 484673
rect 582470 484599 582526 484608
rect 582380 305720 582432 305726
rect 582380 305662 582432 305668
rect 582484 305658 582512 484599
rect 582472 305652 582524 305658
rect 582472 305594 582524 305600
rect 580724 304292 580776 304298
rect 580724 304234 580776 304240
rect 536104 303204 536156 303210
rect 536104 303146 536156 303152
rect 533344 303136 533396 303142
rect 533344 303078 533396 303084
rect 530584 303068 530636 303074
rect 530584 303010 530636 303016
rect 530124 291168 530176 291174
rect 530124 291110 530176 291116
rect 528836 153128 528888 153134
rect 528836 153070 528888 153076
rect 526444 126948 526496 126954
rect 526444 126890 526496 126896
rect 525800 94716 525852 94722
rect 525800 94658 525852 94664
rect 525064 20664 525116 20670
rect 525064 20606 525116 20612
rect 525812 16574 525840 94658
rect 529204 89140 529256 89146
rect 529204 89082 529256 89088
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523040 3596 523092 3602
rect 523040 3538 523092 3544
rect 522304 2984 522356 2990
rect 522304 2926 522356 2932
rect 523052 480 523080 3538
rect 524236 2984 524288 2990
rect 524236 2926 524288 2932
rect 524248 480 524276 2926
rect 525444 480 525472 16546
rect 526180 490 526208 16546
rect 529020 4888 529072 4894
rect 529020 4830 529072 4836
rect 527824 3664 527876 3670
rect 527824 3606 527876 3612
rect 526456 598 526668 626
rect 526456 490 526484 598
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 462 526484 490
rect 526640 480 526668 598
rect 527836 480 527864 3606
rect 529032 480 529060 4830
rect 529216 3058 529244 89082
rect 530596 60722 530624 303010
rect 533356 100706 533384 303078
rect 536116 179382 536144 303146
rect 582472 300960 582524 300966
rect 582472 300902 582524 300908
rect 582380 300892 582432 300898
rect 582380 300834 582432 300840
rect 580172 299532 580224 299538
rect 580172 299474 580224 299480
rect 580184 298761 580212 299474
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580356 298308 580408 298314
rect 580356 298250 580408 298256
rect 580264 298172 580316 298178
rect 580264 298114 580316 298120
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580276 232393 580304 298114
rect 580368 258913 580396 298250
rect 580448 298240 580500 298246
rect 580448 298182 580500 298188
rect 580460 272241 580488 298182
rect 580446 272232 580502 272241
rect 580446 272167 580502 272176
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 206848 580224 206854
rect 580172 206790 580224 206796
rect 580184 205737 580212 206790
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 536104 179376 536156 179382
rect 536104 179318 536156 179324
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 533344 100700 533396 100706
rect 533344 100642 533396 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 550640 98728 550692 98734
rect 550640 98670 550692 98676
rect 532698 95976 532754 95985
rect 532698 95911 532754 95920
rect 530584 60716 530636 60722
rect 530584 60658 530636 60664
rect 530676 60036 530728 60042
rect 530676 59978 530728 59984
rect 530124 3868 530176 3874
rect 530124 3810 530176 3816
rect 529204 3052 529256 3058
rect 529204 2994 529256 3000
rect 530136 480 530164 3810
rect 530688 2990 530716 59978
rect 532712 16574 532740 95911
rect 547142 95840 547198 95849
rect 547142 95775 547198 95784
rect 536840 94648 536892 94654
rect 536840 94590 536892 94596
rect 536104 87848 536156 87854
rect 536104 87790 536156 87796
rect 535460 86284 535512 86290
rect 535460 86226 535512 86232
rect 535472 16574 535500 86226
rect 532712 16546 533752 16574
rect 535472 16546 536052 16574
rect 531320 3052 531372 3058
rect 531320 2994 531372 3000
rect 530676 2984 530728 2990
rect 530676 2926 530728 2932
rect 531332 480 531360 2994
rect 532516 2984 532568 2990
rect 532516 2926 532568 2932
rect 532528 480 532556 2926
rect 533724 480 533752 16546
rect 534908 3528 534960 3534
rect 534908 3470 534960 3476
rect 534920 480 534948 3470
rect 536024 3346 536052 16546
rect 536116 3534 536144 87790
rect 536852 16574 536880 94590
rect 543740 94580 543792 94586
rect 543740 94522 543792 94528
rect 540244 90364 540296 90370
rect 540244 90306 540296 90312
rect 538220 89072 538272 89078
rect 538220 89014 538272 89020
rect 538232 16574 538260 89014
rect 539692 83564 539744 83570
rect 539692 83506 539744 83512
rect 536852 16546 537248 16574
rect 538232 16546 538444 16574
rect 536104 3528 536156 3534
rect 536104 3470 536156 3476
rect 536024 3318 536144 3346
rect 536116 480 536144 3318
rect 537220 480 537248 16546
rect 538416 480 538444 16546
rect 539704 6914 539732 83506
rect 539612 6886 539732 6914
rect 539612 480 539640 6886
rect 540256 3602 540284 90306
rect 543004 87780 543056 87786
rect 543004 87722 543056 87728
rect 540796 3732 540848 3738
rect 540796 3674 540848 3680
rect 540244 3596 540296 3602
rect 540244 3538 540296 3544
rect 540808 480 540836 3674
rect 541992 3596 542044 3602
rect 541992 3538 542044 3544
rect 542004 480 542032 3538
rect 543016 3126 543044 87722
rect 543752 16574 543780 94522
rect 546500 21412 546552 21418
rect 546500 21354 546552 21360
rect 546512 16574 546540 21354
rect 543752 16546 544424 16574
rect 546512 16546 546724 16574
rect 543188 6180 543240 6186
rect 543188 6122 543240 6128
rect 543004 3120 543056 3126
rect 543004 3062 543056 3068
rect 543200 480 543228 6122
rect 544396 480 544424 16546
rect 545488 3120 545540 3126
rect 545488 3062 545540 3068
rect 545500 480 545528 3062
rect 546696 480 546724 16546
rect 547156 3602 547184 95775
rect 547972 87712 548024 87718
rect 547972 87654 548024 87660
rect 547984 16574 548012 87654
rect 550652 16574 550680 98670
rect 554780 98660 554832 98666
rect 554780 98602 554832 98608
rect 554044 93356 554096 93362
rect 554044 93298 554096 93304
rect 553400 84856 553452 84862
rect 553400 84798 553452 84804
rect 553412 16574 553440 84798
rect 547984 16546 548656 16574
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 547144 3596 547196 3602
rect 547144 3538 547196 3544
rect 547880 3460 547932 3466
rect 547880 3402 547932 3408
rect 547892 480 547920 3402
rect 548628 490 548656 16546
rect 550272 3528 550324 3534
rect 550272 3470 550324 3476
rect 548904 598 549116 626
rect 548904 490 548932 598
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 462 548932 490
rect 549088 480 549116 598
rect 550284 480 550312 3470
rect 551020 490 551048 16546
rect 552664 3596 552716 3602
rect 552664 3538 552716 3544
rect 551296 598 551508 626
rect 551296 490 551324 598
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 462 551324 490
rect 551480 480 551508 598
rect 552676 480 552704 3538
rect 553780 480 553808 16546
rect 554056 3126 554084 93298
rect 554792 16574 554820 98602
rect 580262 97200 580318 97209
rect 580262 97135 580318 97144
rect 558184 94512 558236 94518
rect 558184 94454 558236 94460
rect 556252 83496 556304 83502
rect 556252 83438 556304 83444
rect 556264 16574 556292 83438
rect 554792 16546 555004 16574
rect 556264 16546 556936 16574
rect 554044 3120 554096 3126
rect 554044 3062 554096 3068
rect 554976 480 555004 16546
rect 556160 3120 556212 3126
rect 556160 3062 556212 3068
rect 556172 480 556200 3062
rect 556908 490 556936 16546
rect 558196 3466 558224 94454
rect 561680 93288 561732 93294
rect 561680 93230 561732 93236
rect 561692 16574 561720 93230
rect 568580 93220 568632 93226
rect 568580 93162 568632 93168
rect 565820 87644 565872 87650
rect 565820 87586 565872 87592
rect 565084 82204 565136 82210
rect 565084 82146 565136 82152
rect 561692 16546 562088 16574
rect 560392 14680 560444 14686
rect 560392 14622 560444 14628
rect 559288 10532 559340 10538
rect 559288 10474 559340 10480
rect 558552 4820 558604 4826
rect 558552 4762 558604 4768
rect 558184 3460 558236 3466
rect 558184 3402 558236 3408
rect 557184 598 557396 626
rect 557184 490 557212 598
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 462 557212 490
rect 557368 480 557396 598
rect 558564 480 558592 4762
rect 559300 490 559328 10474
rect 559576 598 559788 626
rect 559576 490 559604 598
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559300 462 559604 490
rect 559760 480 559788 598
rect 560404 490 560432 14622
rect 560680 598 560892 626
rect 560680 490 560708 598
rect 559718 -960 559830 480
rect 560404 462 560708 490
rect 560864 480 560892 598
rect 562060 480 562088 16546
rect 564440 14612 564492 14618
rect 564440 14554 564492 14560
rect 563244 10464 563296 10470
rect 563244 10406 563296 10412
rect 563256 480 563284 10406
rect 564452 480 564480 14554
rect 565096 4146 565124 82146
rect 565832 16574 565860 87586
rect 568592 16574 568620 93162
rect 572720 93152 572772 93158
rect 572720 93094 572772 93100
rect 569960 89004 570012 89010
rect 569960 88946 570012 88952
rect 569972 16574 570000 88946
rect 571340 22772 571392 22778
rect 571340 22714 571392 22720
rect 571352 16574 571380 22714
rect 565832 16546 566872 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 571352 16546 571564 16574
rect 565084 4140 565136 4146
rect 565084 4082 565136 4088
rect 565636 3460 565688 3466
rect 565636 3402 565688 3408
rect 565648 480 565676 3402
rect 566844 480 566872 16546
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 568040 480 568068 4082
rect 568684 490 568712 16546
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 16546
rect 571536 480 571564 16546
rect 572732 480 572760 93094
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 575480 80708 575532 80714
rect 575480 80650 575532 80656
rect 575492 16574 575520 80650
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 575492 16546 575888 16574
rect 575112 14544 575164 14550
rect 575112 14486 575164 14492
rect 573456 10396 573508 10402
rect 573456 10338 573508 10344
rect 573468 490 573496 10338
rect 573744 598 573956 626
rect 573744 490 573772 598
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 462 573772 490
rect 573928 480 573956 598
rect 575124 480 575152 14486
rect 575860 490 575888 16546
rect 578608 14476 578660 14482
rect 578608 14418 578660 14424
rect 576952 10328 577004 10334
rect 576952 10270 577004 10276
rect 576136 598 576348 626
rect 576136 490 576164 598
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 462 576164 490
rect 576320 480 576348 598
rect 576964 490 576992 10270
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 576278 -960 576390 480
rect 576964 462 577268 490
rect 577424 480 577452 598
rect 578620 480 578648 14418
rect 580276 3330 580304 97135
rect 582392 6633 582420 300834
rect 582484 46345 582512 300902
rect 582564 82136 582616 82142
rect 582564 82078 582616 82084
rect 582470 46336 582526 46345
rect 582470 46271 582526 46280
rect 582576 16574 582604 82078
rect 582576 16546 583432 16574
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 582196 5024 582248 5030
rect 582196 4966 582248 4972
rect 580264 3324 580316 3330
rect 580264 3266 580316 3272
rect 581000 3324 581052 3330
rect 581000 3266 581052 3272
rect 581012 480 581040 3266
rect 582208 480 582236 4966
rect 583404 480 583432 16546
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 2962 267144 3018 267200
rect 3882 293120 3938 293176
rect 3514 254088 3570 254144
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 2778 97552 2834 97608
rect 12346 94424 12402 94480
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 39302 97144 39358 97200
rect 198462 298832 198518 298888
rect 198554 296792 198610 296848
rect 198462 294616 198518 294672
rect 198646 292576 198702 292632
rect 197358 290400 197414 290456
rect 198554 288360 198610 288416
rect 171138 179188 171140 179208
rect 171140 179188 171192 179208
rect 171192 179188 171194 179208
rect 171138 179152 171194 179188
rect 171782 170448 171838 170504
rect 171874 168136 171930 168192
rect 171966 164464 172022 164520
rect 172426 189896 172482 189952
rect 172426 188672 172482 188728
rect 172426 187312 172482 187368
rect 172426 186088 172482 186144
rect 172426 184764 172428 184784
rect 172428 184764 172480 184784
rect 172480 184764 172482 184784
rect 172426 184728 172482 184764
rect 172334 184320 172390 184376
rect 172426 182960 172482 183016
rect 172426 181736 172482 181792
rect 172426 180512 172482 180568
rect 172426 177948 172482 177984
rect 172426 177928 172428 177948
rect 172428 177928 172480 177948
rect 172480 177928 172482 177948
rect 172242 177384 172298 177440
rect 172242 176024 172298 176080
rect 172426 174800 172482 174856
rect 172426 173576 172482 173632
rect 172426 172388 172428 172408
rect 172428 172388 172480 172408
rect 172480 172388 172482 172408
rect 172426 172352 172482 172388
rect 172426 171028 172428 171048
rect 172428 171028 172480 171048
rect 172480 171028 172482 171048
rect 172426 170992 172482 171028
rect 172242 169088 172298 169144
rect 172426 166640 172482 166696
rect 172058 164056 172114 164112
rect 171690 151544 171746 151600
rect 171506 151000 171562 151056
rect 171598 150456 171654 150512
rect 171690 149912 171746 149968
rect 171690 149404 171692 149424
rect 171692 149404 171744 149424
rect 171744 149404 171746 149424
rect 171690 149368 171746 149404
rect 171690 148280 171746 148336
rect 171506 147736 171562 147792
rect 171506 146648 171562 146704
rect 171506 145016 171562 145072
rect 171414 141924 171416 141944
rect 171416 141924 171468 141944
rect 171468 141924 171470 141944
rect 171414 141888 171470 141924
rect 172242 163512 172298 163568
rect 172150 162288 172206 162344
rect 172426 160928 172482 160984
rect 171782 144064 171838 144120
rect 172334 153720 172390 153776
rect 172242 153176 172298 153232
rect 172426 152632 172482 152688
rect 172334 152088 172390 152144
rect 172242 148860 172244 148880
rect 172244 148860 172296 148880
rect 172296 148860 172298 148880
rect 172242 148824 172298 148860
rect 172426 147192 172482 147248
rect 172334 146140 172336 146160
rect 172336 146140 172388 146160
rect 172388 146140 172390 146160
rect 172334 146104 172390 146140
rect 172426 145560 172482 145616
rect 172426 144472 172482 144528
rect 171966 143520 172022 143576
rect 172242 142976 172298 143032
rect 171598 142432 171654 142488
rect 171506 141344 171562 141400
rect 172426 140800 172482 140856
rect 171506 140256 171562 140312
rect 171690 139748 171692 139768
rect 171692 139748 171744 139768
rect 171744 139748 171746 139768
rect 171690 139712 171746 139748
rect 171874 138624 171930 138680
rect 171690 138080 171746 138136
rect 172426 139168 172482 139224
rect 172426 137536 172482 137592
rect 172242 136992 172298 137048
rect 172334 136448 172390 136504
rect 172426 135904 172482 135960
rect 172242 135360 172298 135416
rect 172242 134816 172298 134872
rect 171874 134272 171930 134328
rect 171690 133864 171746 133920
rect 172518 133320 172574 133376
rect 172426 132776 172482 132832
rect 171138 132232 171194 132288
rect 172426 131688 172482 131744
rect 172334 131144 172390 131200
rect 171322 130600 171378 130656
rect 172242 130056 172298 130112
rect 172150 128968 172206 129024
rect 171966 128424 172022 128480
rect 171782 127336 171838 127392
rect 171506 125160 171562 125216
rect 171874 124616 171930 124672
rect 172058 127880 172114 127936
rect 172426 129512 172482 129568
rect 172334 126792 172390 126848
rect 172242 125740 172244 125760
rect 172244 125740 172296 125760
rect 172296 125740 172298 125760
rect 172242 125704 172298 125740
rect 172426 126248 172482 126304
rect 172150 124228 172206 124264
rect 172150 124208 172152 124228
rect 172152 124208 172204 124228
rect 172204 124208 172206 124228
rect 198186 286184 198242 286240
rect 197358 284144 197414 284200
rect 197910 281968 197966 282024
rect 197542 279928 197598 279984
rect 197358 277752 197414 277808
rect 197542 275712 197598 275768
rect 197358 273536 197414 273592
rect 197542 271496 197598 271552
rect 197634 267280 197690 267336
rect 197358 265104 197414 265160
rect 197358 263064 197414 263120
rect 197358 260908 197414 260944
rect 197358 260888 197360 260908
rect 197360 260888 197412 260908
rect 197412 260888 197414 260908
rect 197358 258848 197414 258904
rect 198002 254632 198058 254688
rect 197910 252456 197966 252512
rect 198094 250416 198150 250472
rect 197542 248240 197598 248296
rect 198094 246200 198150 246256
rect 197542 244024 197598 244080
rect 197542 239808 197598 239864
rect 197542 235592 197598 235648
rect 197358 233552 197414 233608
rect 197358 229336 197414 229392
rect 197542 227296 197598 227352
rect 197358 225120 197414 225176
rect 198002 223080 198058 223136
rect 197358 220924 197414 220960
rect 197358 220904 197360 220924
rect 197360 220904 197412 220924
rect 197412 220904 197414 220924
rect 197542 218864 197598 218920
rect 197358 216708 197414 216744
rect 197358 216688 197360 216708
rect 197360 216688 197412 216708
rect 197412 216688 197414 216708
rect 197358 214648 197414 214704
rect 197358 212472 197414 212528
rect 197358 210432 197414 210488
rect 197358 208256 197414 208312
rect 197358 206216 197414 206272
rect 197358 202000 197414 202056
rect 197542 199824 197598 199880
rect 197358 197784 197414 197840
rect 197542 195608 197598 195664
rect 197358 193568 197414 193624
rect 197358 189352 197414 189408
rect 197358 187176 197414 187232
rect 197358 182960 197414 183016
rect 197358 178744 197414 178800
rect 197358 176724 197414 176760
rect 197358 176704 197360 176724
rect 197360 176704 197412 176724
rect 197412 176704 197414 176724
rect 197726 174528 197782 174584
rect 197358 172524 197360 172544
rect 197360 172524 197412 172544
rect 197412 172524 197414 172544
rect 197358 172488 197414 172524
rect 197450 170312 197506 170368
rect 197358 168272 197414 168328
rect 197542 164056 197598 164112
rect 197542 159840 197598 159896
rect 197358 157800 197414 157856
rect 197542 155624 197598 155680
rect 197358 153584 197414 153640
rect 197542 151408 197598 151464
rect 197358 149368 197414 149424
rect 197634 147192 197690 147248
rect 197358 145152 197414 145208
rect 197358 142976 197414 143032
rect 197358 140936 197414 140992
rect 197358 138760 197414 138816
rect 197358 136720 197414 136776
rect 198462 269340 198518 269376
rect 198462 269320 198464 269340
rect 198464 269320 198516 269340
rect 198516 269320 198518 269340
rect 198370 256708 198372 256728
rect 198372 256708 198424 256728
rect 198424 256708 198426 256728
rect 198370 256672 198426 256708
rect 198278 241984 198334 242040
rect 198462 237788 198518 237824
rect 198462 237768 198464 237788
rect 198464 237768 198516 237788
rect 198516 237768 198518 237788
rect 198738 231512 198794 231568
rect 198278 204040 198334 204096
rect 198278 191392 198334 191448
rect 198462 185136 198518 185192
rect 198278 180940 198334 180976
rect 198278 180920 198280 180940
rect 198280 180920 198332 180940
rect 198332 180920 198334 180940
rect 198462 166232 198518 166288
rect 213826 299376 213882 299432
rect 214378 299240 214434 299296
rect 216034 299376 216090 299432
rect 216954 299376 217010 299432
rect 214562 299276 214564 299296
rect 214564 299276 214616 299296
rect 214616 299276 214618 299296
rect 214562 299240 214618 299276
rect 224406 299276 224408 299296
rect 224408 299276 224460 299296
rect 224460 299276 224462 299296
rect 224406 299240 224462 299276
rect 302882 298424 302938 298480
rect 302790 295332 302792 295352
rect 302792 295332 302844 295352
rect 302844 295332 302846 295352
rect 302790 295296 302846 295332
rect 302238 289212 302240 289232
rect 302240 289212 302292 289232
rect 302292 289212 302294 289232
rect 302238 289176 302294 289212
rect 302238 286048 302294 286104
rect 302790 283056 302846 283112
rect 302422 279928 302478 279984
rect 302790 276800 302846 276856
rect 302698 273808 302754 273864
rect 302974 292304 303030 292360
rect 303066 270680 303122 270736
rect 302882 267688 302938 267744
rect 302698 264560 302754 264616
rect 302330 261432 302386 261488
rect 302606 258440 302662 258496
rect 302790 255312 302846 255368
rect 302790 249192 302846 249248
rect 302514 246064 302570 246120
rect 302974 252184 303030 252240
rect 303250 252184 303306 252240
rect 303250 243072 303306 243128
rect 302882 239944 302938 240000
rect 302790 236816 302846 236872
rect 302698 233824 302754 233880
rect 302790 230696 302846 230752
rect 302790 227568 302846 227624
rect 302330 224576 302386 224632
rect 302330 221448 302386 221504
rect 302422 218320 302478 218376
rect 302882 212200 302938 212256
rect 302238 206116 302240 206136
rect 302240 206116 302292 206136
rect 302292 206116 302294 206136
rect 302238 206080 302294 206116
rect 302790 196832 302846 196888
rect 302606 193704 302662 193760
rect 302422 190712 302478 190768
rect 302790 184592 302846 184648
rect 302698 181464 302754 181520
rect 302238 175344 302294 175400
rect 302790 169088 302846 169144
rect 302790 166096 302846 166152
rect 302790 162968 302846 163024
rect 198094 162016 198150 162072
rect 302514 159840 302570 159896
rect 303066 215328 303122 215384
rect 303066 209208 303122 209264
rect 302974 202952 303030 203008
rect 302790 156848 302846 156904
rect 303434 199960 303490 200016
rect 303066 187584 303122 187640
rect 303342 178336 303398 178392
rect 303066 172216 303122 172272
rect 302790 153720 302846 153776
rect 302790 150728 302846 150784
rect 302698 147600 302754 147656
rect 302790 144472 302846 144528
rect 302330 141480 302386 141536
rect 302882 138352 302938 138408
rect 197726 134544 197782 134600
rect 197358 132524 197414 132560
rect 197358 132504 197360 132524
rect 197360 132504 197412 132524
rect 197412 132504 197414 132524
rect 302514 132232 302570 132288
rect 197358 130328 197414 130384
rect 197358 128308 197414 128344
rect 197358 128288 197360 128308
rect 197360 128288 197412 128308
rect 197412 128288 197414 128308
rect 197634 126112 197690 126168
rect 302422 126112 302478 126168
rect 302698 129104 302754 129160
rect 302974 135224 303030 135280
rect 197358 124108 197360 124128
rect 197360 124108 197412 124128
rect 197412 124108 197414 124128
rect 197358 124072 197414 124108
rect 302238 122984 302294 123040
rect 197450 121896 197506 121952
rect 197358 119856 197414 119912
rect 197634 117680 197690 117736
rect 198554 115640 198610 115696
rect 197542 113464 197598 113520
rect 197358 111424 197414 111480
rect 197542 109248 197598 109304
rect 198002 107208 198058 107264
rect 197450 105032 197506 105088
rect 198002 102992 198058 103048
rect 198002 100952 198058 101008
rect 195334 97824 195390 97880
rect 200854 97824 200910 97880
rect 202050 94424 202106 94480
rect 203430 97144 203486 97200
rect 280158 97280 280214 97336
rect 281998 97588 282000 97608
rect 282000 97588 282052 97608
rect 282052 97588 282054 97608
rect 281998 97552 282054 97588
rect 285862 97552 285918 97608
rect 289910 95920 289966 95976
rect 293130 95784 293186 95840
rect 297086 96600 297142 96656
rect 297914 97416 297970 97472
rect 297730 97144 297786 97200
rect 302514 119856 302570 119912
rect 302606 116864 302662 116920
rect 302514 110608 302570 110664
rect 302790 107616 302846 107672
rect 302974 113736 303030 113792
rect 302882 104488 302938 104544
rect 302790 101496 302846 101552
rect 298742 96600 298798 96656
rect 371238 585656 371294 585712
rect 371698 585112 371754 585168
rect 371422 584568 371478 584624
rect 371330 581848 371386 581904
rect 371790 582392 371846 582448
rect 372158 582392 372214 582448
rect 371606 581304 371662 581360
rect 371698 580760 371754 580816
rect 371514 580216 371570 580272
rect 371330 578584 371386 578640
rect 369858 569200 369914 569256
rect 369306 568656 369362 568712
rect 362866 553424 362922 553480
rect 364890 553424 364946 553480
rect 369306 566480 369362 566536
rect 369398 511828 369454 511864
rect 369398 511808 369400 511828
rect 369400 511808 369452 511828
rect 369452 511808 369454 511828
rect 369950 567160 370006 567216
rect 369858 512896 369914 512952
rect 369490 507456 369546 507512
rect 365166 484064 365222 484120
rect 362866 482160 362922 482216
rect 369766 488144 369822 488200
rect 369306 423136 369362 423192
rect 369306 420960 369362 421016
rect 369490 425176 369546 425232
rect 369398 413888 369454 413944
rect 362774 411984 362830 412040
rect 365166 411984 365222 412040
rect 362498 340448 362554 340504
rect 365166 340448 365222 340504
rect 370134 564168 370190 564224
rect 369950 509360 370006 509416
rect 369858 425856 369914 425912
rect 370042 504872 370098 504928
rect 369950 423544 370006 423600
rect 370226 561992 370282 562048
rect 370134 501880 370190 501936
rect 370042 421640 370098 421696
rect 369950 417696 370006 417752
rect 369858 411576 369914 411632
rect 356702 266056 356758 266112
rect 358174 266192 358230 266248
rect 369306 359760 369362 359816
rect 369766 358808 369822 358864
rect 370318 561448 370374 561504
rect 370226 497256 370282 497312
rect 370134 420144 370190 420200
rect 370042 360848 370098 360904
rect 369950 353504 370006 353560
rect 369858 340856 369914 340912
rect 369398 297492 369454 297528
rect 369398 297472 369400 297492
rect 369400 297472 369452 297492
rect 369452 297472 369454 297492
rect 369858 297372 369860 297392
rect 369860 297372 369912 297392
rect 369912 297372 369914 297392
rect 369858 297336 369914 297372
rect 369398 295840 369454 295896
rect 369858 295860 369914 295896
rect 369858 295840 369860 295860
rect 369860 295840 369912 295860
rect 369912 295840 369914 295860
rect 369490 291896 369546 291952
rect 369398 283348 369454 283384
rect 369398 283328 369400 283348
rect 369400 283328 369452 283348
rect 369452 283328 369454 283348
rect 369398 280744 369454 280800
rect 362866 266192 362922 266248
rect 364890 265784 364946 265840
rect 367834 225684 367890 225720
rect 367834 225664 367836 225684
rect 367836 225664 367888 225684
rect 367888 225664 367890 225684
rect 369950 287816 370006 287872
rect 369858 284416 369914 284472
rect 369674 277480 369730 277536
rect 369398 224168 369454 224224
rect 369490 223624 369546 223680
rect 365166 196424 365222 196480
rect 362866 194520 362922 194576
rect 370410 558184 370466 558240
rect 370318 496168 370374 496224
rect 370502 556144 370558 556200
rect 370410 489232 370466 489288
rect 370962 511164 370964 511184
rect 370964 511164 371016 511184
rect 371016 511164 371018 511184
rect 370962 511128 371018 511164
rect 370962 510060 371018 510096
rect 370962 510040 370964 510060
rect 370964 510040 371016 510060
rect 371016 510040 371018 510060
rect 370962 506524 371018 506560
rect 370962 506504 370964 506524
rect 370964 506504 371016 506524
rect 371016 506504 371018 506524
rect 370962 504212 371018 504248
rect 370962 504192 370964 504212
rect 370964 504192 371016 504212
rect 371016 504192 371018 504212
rect 370962 503140 370964 503160
rect 370964 503140 371016 503160
rect 371016 503140 371018 503160
rect 370962 503104 371018 503140
rect 370962 499604 370964 499624
rect 370964 499604 371016 499624
rect 371016 499604 371018 499624
rect 370962 499568 371018 499604
rect 370962 498500 371018 498536
rect 370962 498480 370964 498500
rect 370964 498480 371016 498500
rect 371016 498480 371018 498500
rect 370686 496168 370742 496224
rect 370962 494944 371018 495000
rect 370962 493856 371018 493912
rect 370778 492632 370834 492688
rect 370502 484608 370558 484664
rect 370410 422456 370466 422512
rect 370226 417968 370282 418024
rect 370226 414160 370282 414216
rect 370134 357856 370190 357912
rect 370042 278024 370098 278080
rect 370318 367104 370374 367160
rect 370870 491544 370926 491600
rect 370962 490340 371018 490376
rect 370962 490320 370964 490340
rect 370964 490320 371016 490340
rect 371016 490320 371018 490340
rect 370962 485696 371018 485752
rect 371146 482876 371148 482896
rect 371148 482876 371200 482896
rect 371200 482876 371202 482896
rect 371146 482840 371202 482876
rect 371422 577496 371478 577552
rect 371606 579708 371608 579728
rect 371608 579708 371660 579728
rect 371660 579708 371662 579728
rect 371606 579672 371662 579708
rect 371698 579128 371754 579184
rect 371698 578040 371754 578096
rect 371606 576972 371662 577008
rect 371606 576952 371608 576972
rect 371608 576952 371660 576972
rect 371660 576952 371662 576972
rect 371330 441768 371386 441824
rect 371238 441088 371294 441144
rect 371238 440408 371294 440464
rect 371698 576408 371754 576464
rect 371882 576000 371938 576056
rect 371606 575456 371662 575512
rect 371790 574912 371846 574968
rect 371606 571648 371662 571704
rect 371698 571104 371754 571160
rect 371514 570560 371570 570616
rect 371606 570036 371662 570072
rect 371606 570016 371608 570036
rect 371608 570016 371660 570036
rect 371660 570016 371662 570036
rect 371514 568384 371570 568440
rect 371606 567840 371662 567896
rect 371422 440544 371478 440600
rect 371974 573824 372030 573880
rect 371238 427352 371294 427408
rect 371054 425448 371110 425504
rect 371238 424904 371294 424960
rect 371146 423272 371202 423328
rect 370870 417424 370926 417480
rect 370686 414160 370742 414216
rect 370502 412120 370558 412176
rect 370594 368328 370650 368384
rect 370410 363704 370466 363760
rect 370778 363704 370834 363760
rect 370686 357876 370742 357912
rect 370686 357856 370688 357876
rect 370688 357856 370740 357876
rect 370740 357856 370742 357876
rect 370594 353232 370650 353288
rect 370686 350920 370742 350976
rect 370502 347520 370558 347576
rect 370226 345228 370282 345264
rect 370226 345208 370228 345228
rect 370228 345208 370280 345228
rect 370280 345208 370282 345228
rect 370226 340584 370282 340640
rect 370042 276936 370098 276992
rect 369950 267960 370006 268016
rect 370502 295024 370558 295080
rect 370410 285368 370466 285424
rect 370318 278840 370374 278896
rect 370594 294480 370650 294536
rect 370686 292848 370742 292904
rect 371238 415248 371294 415304
rect 371238 413616 371294 413672
rect 370962 369416 371018 369472
rect 371606 437824 371662 437880
rect 371790 566228 371846 566264
rect 371790 566208 371792 566228
rect 371792 566208 371844 566228
rect 371844 566208 371846 566228
rect 371790 565836 371792 565856
rect 371792 565836 371844 565856
rect 371844 565836 371846 565856
rect 371790 565800 371846 565836
rect 371790 564732 371846 564768
rect 371790 564712 371792 564732
rect 371792 564712 371844 564732
rect 371844 564712 371846 564732
rect 371790 563100 371846 563136
rect 371790 563080 371792 563100
rect 371792 563080 371844 563100
rect 371844 563080 371846 563100
rect 371790 562556 371846 562592
rect 371790 562536 371792 562556
rect 371792 562536 371844 562556
rect 371844 562536 371846 562556
rect 371790 560924 371846 560960
rect 371790 560904 371792 560924
rect 371792 560904 371844 560924
rect 371844 560904 371846 560924
rect 371790 560380 371846 560416
rect 371790 560360 371792 560380
rect 371792 560360 371844 560380
rect 371844 560360 371846 560380
rect 371882 559816 371938 559872
rect 371790 559272 371846 559328
rect 371790 558728 371846 558784
rect 371790 557640 371846 557696
rect 371790 556552 371846 556608
rect 371882 440408 371938 440464
rect 371790 438368 371846 438424
rect 371698 437280 371754 437336
rect 371606 436736 371662 436792
rect 371790 436192 371846 436248
rect 371606 435648 371662 435704
rect 371698 435104 371754 435160
rect 371606 434580 371662 434616
rect 371606 434560 371608 434580
rect 371608 434560 371660 434580
rect 371660 434560 371662 434580
rect 371698 434016 371754 434072
rect 371790 433472 371846 433528
rect 371698 432928 371754 432984
rect 371606 432384 371662 432440
rect 371606 431976 371662 432032
rect 371514 430888 371570 430944
rect 370962 366016 371018 366072
rect 370962 364812 371018 364848
rect 370962 364792 370964 364812
rect 370964 364792 371016 364812
rect 371016 364792 371018 364812
rect 370962 362500 371018 362536
rect 370962 362480 370964 362500
rect 370964 362480 371016 362500
rect 371016 362480 371018 362500
rect 370962 356788 371018 356824
rect 370962 356768 370964 356788
rect 370964 356768 371016 356788
rect 371016 356768 371018 356788
rect 370962 355564 371018 355600
rect 370962 355544 370964 355564
rect 370964 355544 371016 355564
rect 371016 355544 371018 355564
rect 370962 354476 371018 354512
rect 370962 354456 370964 354476
rect 370964 354456 371016 354476
rect 371016 354456 371018 354476
rect 370870 352164 370926 352200
rect 370870 352144 370872 352164
rect 370872 352144 370924 352164
rect 370924 352144 370926 352164
rect 370962 349852 371018 349888
rect 370962 349832 370964 349852
rect 370964 349832 371016 349852
rect 371016 349832 371018 349852
rect 370962 348644 370964 348664
rect 370964 348644 371016 348664
rect 371016 348644 371018 348664
rect 370962 348608 371018 348644
rect 370962 346316 371018 346352
rect 370962 346296 370964 346316
rect 370964 346296 371016 346316
rect 371016 346296 371018 346316
rect 370962 344004 371018 344040
rect 370962 343984 370964 344004
rect 370964 343984 371016 344004
rect 371016 343984 371018 344004
rect 370962 342916 371018 342952
rect 370962 342896 370964 342916
rect 370964 342896 371016 342916
rect 371016 342896 371018 342916
rect 371238 298016 371294 298072
rect 371330 297744 371386 297800
rect 371422 296656 371478 296712
rect 371422 295296 371478 295352
rect 371330 294480 371386 294536
rect 371330 293392 371386 293448
rect 371238 292848 371294 292904
rect 371238 292304 371294 292360
rect 371238 289584 371294 289640
rect 371330 287544 371386 287600
rect 371698 431432 371754 431488
rect 371698 430616 371754 430672
rect 371606 427100 371662 427136
rect 371606 427080 371608 427100
rect 371608 427080 371660 427100
rect 371660 427080 371662 427100
rect 371606 426572 371608 426592
rect 371608 426572 371660 426592
rect 371660 426572 371662 426592
rect 371606 426536 371662 426572
rect 371606 426028 371608 426048
rect 371608 426028 371660 426048
rect 371660 426028 371662 426048
rect 371606 425992 371662 426028
rect 371606 423836 371662 423872
rect 371606 423816 371608 423836
rect 371608 423816 371660 423836
rect 371660 423816 371662 423836
rect 370778 278840 370834 278896
rect 370318 219680 370374 219736
rect 370318 218476 370374 218512
rect 370318 218456 370320 218476
rect 370320 218456 370372 218476
rect 370372 218456 370374 218476
rect 370134 215056 370190 215112
rect 369950 196832 370006 196888
rect 369306 151680 369362 151736
rect 369490 151272 369546 151328
rect 369582 150728 369638 150784
rect 369398 143792 369454 143848
rect 369306 136584 369362 136640
rect 369306 134952 369362 135008
rect 371514 287000 371570 287056
rect 371882 430616 371938 430672
rect 371790 297200 371846 297256
rect 371698 293936 371754 293992
rect 371698 291796 371700 291816
rect 371700 291796 371752 291816
rect 371752 291796 371754 291816
rect 371698 291760 371754 291796
rect 371698 291236 371754 291272
rect 371698 291216 371700 291236
rect 371700 291216 371752 291236
rect 371752 291216 371754 291236
rect 371698 290672 371754 290728
rect 372066 573280 372122 573336
rect 371974 429800 372030 429856
rect 372434 574368 372490 574424
rect 372250 572736 372306 572792
rect 372250 556008 372306 556064
rect 372158 430344 372214 430400
rect 372066 429256 372122 429312
rect 372526 565256 372582 565312
rect 372710 563624 372766 563680
rect 372526 500792 372582 500848
rect 372802 557096 372858 557152
rect 372526 486920 372582 486976
rect 372250 428712 372306 428768
rect 371974 422184 372030 422240
rect 371974 420724 371976 420744
rect 371976 420724 372028 420744
rect 372028 420724 372030 420744
rect 371974 420688 372030 420724
rect 371974 419092 371976 419112
rect 371976 419092 372028 419112
rect 372028 419092 372030 419112
rect 371974 419056 372030 419092
rect 371974 416880 372030 416936
rect 371974 416372 371976 416392
rect 371976 416372 372028 416392
rect 372028 416372 372030 416392
rect 371974 416336 372030 416372
rect 371974 415792 372030 415848
rect 371974 414740 371976 414760
rect 371976 414740 372028 414760
rect 372028 414740 372030 414760
rect 371974 414704 372030 414740
rect 372434 419600 372490 419656
rect 372158 418512 372214 418568
rect 371790 290128 371846 290184
rect 371698 289040 371754 289096
rect 371698 288532 371700 288552
rect 371700 288532 371752 288552
rect 371752 288532 371754 288552
rect 371698 288496 371754 288532
rect 371882 288088 371938 288144
rect 372066 412548 372122 412584
rect 372066 412528 372068 412548
rect 372068 412528 372120 412548
rect 372120 412528 372122 412548
rect 372250 298016 372306 298072
rect 372066 295296 372122 295352
rect 372158 295024 372214 295080
rect 372342 296132 372398 296168
rect 372342 296112 372344 296132
rect 372344 296112 372396 296132
rect 372396 296112 372398 296132
rect 372618 424360 372674 424416
rect 372802 413072 372858 413128
rect 371974 286456 372030 286512
rect 371146 285912 371202 285968
rect 372342 285368 372398 285424
rect 372434 284824 372490 284880
rect 372250 284316 372252 284336
rect 372252 284316 372304 284336
rect 372304 284316 372306 284336
rect 372250 284280 372306 284316
rect 371514 283192 371570 283248
rect 371606 282648 371662 282704
rect 371698 282104 371754 282160
rect 371238 281560 371294 281616
rect 371514 281560 371570 281616
rect 371514 281016 371570 281072
rect 371238 225664 371294 225720
rect 371422 279928 371478 279984
rect 371606 279404 371662 279440
rect 371606 279384 371608 279404
rect 371608 279384 371660 279404
rect 371660 279384 371662 279404
rect 371606 278316 371662 278352
rect 371606 278296 371608 278316
rect 371608 278296 371660 278316
rect 371660 278296 371662 278316
rect 371422 277344 371478 277400
rect 372434 276276 372490 276312
rect 372434 276256 372436 276276
rect 372436 276256 372488 276276
rect 372488 276256 372490 276276
rect 371606 275748 371608 275768
rect 371608 275748 371660 275768
rect 371660 275748 371662 275768
rect 371606 275712 371662 275748
rect 372158 275204 372160 275224
rect 372160 275204 372212 275224
rect 372212 275204 372214 275224
rect 372158 275168 372214 275204
rect 371514 274080 371570 274136
rect 371606 273572 371608 273592
rect 371608 273572 371660 273592
rect 371660 273572 371662 273592
rect 371606 273536 371662 273572
rect 373078 421232 373134 421288
rect 372802 341672 372858 341728
rect 372986 278024 373042 278080
rect 371698 272992 371754 273048
rect 371882 272448 371938 272504
rect 371790 271904 371846 271960
rect 371422 269184 371478 269240
rect 370962 217388 371018 217424
rect 370962 217368 370964 217388
rect 370964 217368 371016 217388
rect 371016 217368 371018 217388
rect 370962 216180 370964 216200
rect 370964 216180 371016 216200
rect 371016 216180 371018 216200
rect 370962 216144 371018 216180
rect 370686 215076 370742 215112
rect 370686 215056 370688 215076
rect 370688 215056 370740 215076
rect 370740 215056 370742 215076
rect 370962 213852 371018 213888
rect 370962 213832 370964 213852
rect 370964 213832 371016 213852
rect 371016 213832 371018 213852
rect 370962 211556 370964 211576
rect 370964 211556 371016 211576
rect 371016 211556 371018 211576
rect 370962 211520 371018 211556
rect 370962 210432 371018 210488
rect 370962 209228 371018 209264
rect 370962 209208 370964 209228
rect 370964 209208 371016 209228
rect 371016 209208 371018 209228
rect 370962 208140 371018 208176
rect 370962 208120 370964 208140
rect 370964 208120 371016 208140
rect 371016 208120 371018 208140
rect 371238 205808 371294 205864
rect 370962 197668 371018 197704
rect 370962 197648 370964 197668
rect 370964 197648 371016 197668
rect 371016 197648 371018 197668
rect 370870 196560 370926 196616
rect 370410 149912 370466 149968
rect 370318 148824 370374 148880
rect 370226 141888 370282 141944
rect 370594 140800 370650 140856
rect 370502 140256 370558 140312
rect 370134 139712 370190 139768
rect 370042 133592 370098 133648
rect 369858 132368 369914 132424
rect 369490 131960 369546 132016
rect 369398 131416 369454 131472
rect 370042 130192 370098 130248
rect 369858 129104 369914 129160
rect 369306 128560 369362 128616
rect 369398 126384 369454 126440
rect 362774 123936 362830 123992
rect 365166 123936 365222 123992
rect 369950 128560 370006 128616
rect 370318 130056 370374 130112
rect 370226 127880 370282 127936
rect 370134 127336 370190 127392
rect 369858 124344 369914 124400
rect 369950 123936 370006 123992
rect 370410 126248 370466 126304
rect 370502 125704 370558 125760
rect 371330 202272 371386 202328
rect 371238 152904 371294 152960
rect 371238 149368 371294 149424
rect 371790 270816 371846 270872
rect 371974 270272 372030 270328
rect 371882 269728 371938 269784
rect 371514 221992 371570 222048
rect 371790 206896 371846 206952
rect 371514 201184 371570 201240
rect 371422 198872 371478 198928
rect 371330 147736 371386 147792
rect 371330 147228 371332 147248
rect 371332 147228 371384 147248
rect 371384 147228 371386 147248
rect 371330 147192 371386 147228
rect 371330 145596 371332 145616
rect 371332 145596 371384 145616
rect 371384 145596 371386 145616
rect 371330 145560 371386 145596
rect 371330 145016 371386 145072
rect 371330 144508 371332 144528
rect 371332 144508 371384 144528
rect 371384 144508 371386 144528
rect 371330 144472 371386 144508
rect 371330 144100 371332 144120
rect 371332 144100 371384 144120
rect 371384 144100 371386 144120
rect 371330 144064 371386 144100
rect 371330 142432 371386 142488
rect 371330 138080 371386 138136
rect 371330 137572 371332 137592
rect 371332 137572 371384 137592
rect 371384 137572 371386 137592
rect 371330 137536 371386 137572
rect 371238 126384 371294 126440
rect 371606 199960 371662 200016
rect 371514 132776 371570 132832
rect 371698 138624 371754 138680
rect 371698 134308 371700 134328
rect 371700 134308 371752 134328
rect 371752 134308 371754 134328
rect 371698 134272 371754 134308
rect 372526 271360 372582 271416
rect 372802 274624 372858 274680
rect 372526 269864 372582 269920
rect 372526 268640 372582 268696
rect 372526 223080 372582 223136
rect 372342 220768 372398 220824
rect 372250 205808 372306 205864
rect 372250 204584 372306 204640
rect 372158 203496 372214 203552
rect 372066 202272 372122 202328
rect 371974 201184 372030 201240
rect 371790 128968 371846 129024
rect 372434 168952 372490 169008
rect 372802 212744 372858 212800
rect 372158 158752 372214 158808
rect 371974 146648 372030 146704
rect 371974 146104 372030 146160
rect 371974 143012 371976 143032
rect 371976 143012 372028 143032
rect 372028 143012 372030 143032
rect 371974 142976 372030 143012
rect 371974 141344 372030 141400
rect 371974 135904 372030 135960
rect 371882 128560 371938 128616
rect 372158 139168 372214 139224
rect 375102 289856 375158 289912
rect 375194 289448 375250 289504
rect 372342 135360 372398 135416
rect 372526 133864 372582 133920
rect 372802 136992 372858 137048
rect 373998 129512 374054 129568
rect 372066 127880 372122 127936
rect 371698 126384 371754 126440
rect 371606 125704 371662 125760
rect 371422 125160 371478 125216
rect 370870 124208 370926 124264
rect 374734 220768 374790 220824
rect 375102 231784 375158 231840
rect 375194 231648 375250 231704
rect 445666 585384 445722 585440
rect 444746 584296 444802 584352
rect 442998 583072 443054 583128
rect 441618 577088 441674 577144
rect 441618 559408 441674 559464
rect 441802 573280 441858 573336
rect 441710 556844 441766 556880
rect 441710 556824 441712 556844
rect 441712 556824 441764 556844
rect 441764 556824 441766 556844
rect 435178 553424 435234 553480
rect 436742 553424 436798 553480
rect 441710 507320 441766 507376
rect 441618 504600 441674 504656
rect 435178 483928 435234 483984
rect 436742 483928 436798 483984
rect 441066 409536 441122 409592
rect 434902 408584 434958 408640
rect 436834 408584 436890 408640
rect 441894 567568 441950 567624
rect 441802 492496 441858 492552
rect 441986 561720 442042 561776
rect 441894 489640 441950 489696
rect 442078 558864 442134 558920
rect 441986 486920 442042 486976
rect 443090 580760 443146 580816
rect 442998 496440 443054 496496
rect 444746 579692 444802 579728
rect 444746 579672 444748 579692
rect 444748 579672 444800 579692
rect 444800 579672 444802 579692
rect 444930 578468 444986 578504
rect 444930 578448 444932 578468
rect 444932 578448 444984 578468
rect 444984 578448 444986 578468
rect 444746 576136 444802 576192
rect 444562 575048 444618 575104
rect 444838 571532 444894 571568
rect 444838 571512 444840 571532
rect 444840 571512 444892 571532
rect 444892 571512 444894 571532
rect 443182 570424 443238 570480
rect 443090 495352 443146 495408
rect 442906 494808 442962 494864
rect 442078 485152 442134 485208
rect 441802 435512 441858 435568
rect 441342 368872 441398 368928
rect 441618 369416 441674 369472
rect 441342 367820 441344 367840
rect 441344 367820 441396 367840
rect 441396 367820 441398 367840
rect 441342 367784 441398 367820
rect 441618 367784 441674 367840
rect 441710 363976 441766 364032
rect 441618 361256 441674 361312
rect 441894 429256 441950 429312
rect 441710 351056 441766 351112
rect 442078 428712 442134 428768
rect 441986 423952 442042 424008
rect 441894 348472 441950 348528
rect 442998 493856 443054 493912
rect 442538 492224 442594 492280
rect 442446 435648 442502 435704
rect 442630 485696 442686 485752
rect 442538 429800 442594 429856
rect 442354 424088 442410 424144
rect 442262 422864 442318 422920
rect 442078 419464 442134 419520
rect 441986 345752 442042 345808
rect 441894 343576 441950 343632
rect 441802 343032 441858 343088
rect 441618 340892 441620 340912
rect 441620 340892 441672 340912
rect 441672 340892 441674 340912
rect 441618 340856 441674 340892
rect 431866 338000 431922 338056
rect 431774 337864 431830 337920
rect 400126 298152 400182 298208
rect 436558 340040 436614 340096
rect 434856 339904 434912 339960
rect 436558 338000 436614 338056
rect 434810 337864 434866 337920
rect 440790 340040 440846 340096
rect 441710 296928 441766 296984
rect 441710 295976 441766 296032
rect 444930 569200 444986 569256
rect 443274 566888 443330 566944
rect 444470 565800 444526 565856
rect 444378 564596 444434 564632
rect 444378 564576 444380 564596
rect 444380 564576 444432 564596
rect 444432 564576 444434 564596
rect 444378 561196 444434 561232
rect 444378 561176 444380 561196
rect 444380 561176 444432 561196
rect 444432 561176 444434 561196
rect 444378 557660 444434 557696
rect 444378 557640 444380 557660
rect 444380 557640 444432 557660
rect 444432 557640 444434 557660
rect 445666 563488 445722 563544
rect 444378 513748 444380 513768
rect 444380 513748 444432 513768
rect 444432 513748 444434 513768
rect 444378 513712 444434 513748
rect 444838 513168 444894 513224
rect 444378 512624 444434 512680
rect 443182 490592 443238 490648
rect 443826 496440 443882 496496
rect 443642 495352 443698 495408
rect 443550 491680 443606 491736
rect 443458 488960 443514 489016
rect 443274 486376 443330 486432
rect 442998 433336 443054 433392
rect 442170 415928 442226 415984
rect 442630 415928 442686 415984
rect 442078 343304 442134 343360
rect 442262 369164 442318 369200
rect 442262 369144 442264 369164
rect 442264 369144 442316 369164
rect 442316 369144 442318 369164
rect 442262 366968 442318 367024
rect 442170 341400 442226 341456
rect 442446 365880 442502 365936
rect 443090 431060 443092 431080
rect 443092 431060 443144 431080
rect 443144 431060 443146 431080
rect 443090 431024 443146 431060
rect 442998 349832 443054 349888
rect 443366 484744 443422 484800
rect 443274 418240 443330 418296
rect 443918 490048 443974 490104
rect 443826 439048 443882 439104
rect 444562 512080 444618 512136
rect 444194 439068 444250 439104
rect 444194 439048 444196 439068
rect 444196 439048 444248 439068
rect 444248 439048 444250 439068
rect 444378 436756 444434 436792
rect 444378 436736 444380 436756
rect 444380 436736 444432 436756
rect 444432 436736 444434 436756
rect 443550 425176 443606 425232
rect 443918 425176 443974 425232
rect 443458 418240 443514 418296
rect 443366 414840 443422 414896
rect 443366 350512 443422 350568
rect 443090 348744 443146 348800
rect 442998 342760 443054 342816
rect 441986 286456 442042 286512
rect 441802 275712 441858 275768
rect 443090 341400 443146 341456
rect 442998 274352 443054 274408
rect 443826 421776 443882 421832
rect 444194 414860 444250 414896
rect 444194 414840 444196 414860
rect 444196 414840 444248 414860
rect 444248 414840 444250 414860
rect 443550 346024 443606 346080
rect 444470 434444 444526 434480
rect 444470 434424 444472 434444
rect 444472 434424 444524 434444
rect 444524 434424 444526 434444
rect 444470 432112 444526 432168
rect 444470 419484 444526 419520
rect 444470 419464 444472 419484
rect 444472 419464 444524 419484
rect 444524 419464 444526 419484
rect 444378 368600 444434 368656
rect 444286 366424 444342 366480
rect 444194 365336 444250 365392
rect 443734 349832 443790 349888
rect 443642 344392 443698 344448
rect 443458 342760 443514 342816
rect 443366 291760 443422 291816
rect 443642 292848 443698 292904
rect 444746 510448 444802 510504
rect 444654 498616 444710 498672
rect 444654 492768 444710 492824
rect 444654 487892 444710 487928
rect 444654 487872 444656 487892
rect 444656 487872 444708 487892
rect 444708 487872 444710 487892
rect 444654 484220 444710 484256
rect 444654 484200 444656 484220
rect 444656 484200 444708 484220
rect 444708 484200 444710 484220
rect 444654 437980 444710 438016
rect 444654 437960 444656 437980
rect 444656 437960 444708 437980
rect 444708 437960 444710 437980
rect 444654 417172 444710 417208
rect 444654 417152 444656 417172
rect 444656 417152 444708 417172
rect 444708 417152 444710 417172
rect 445666 511536 445722 511592
rect 445390 510992 445446 511048
rect 445298 504056 445354 504112
rect 445114 503512 445170 503568
rect 445022 502968 445078 503024
rect 445206 502424 445262 502480
rect 445298 501336 445354 501392
rect 445114 485732 445116 485752
rect 445116 485732 445168 485752
rect 445168 485732 445170 485752
rect 445114 485696 445170 485732
rect 444930 369688 444986 369744
rect 444838 369144 444894 369200
rect 444654 365880 444710 365936
rect 444930 364792 444986 364848
rect 444470 362616 444526 362672
rect 445298 494264 445354 494320
rect 445298 493348 445300 493368
rect 445300 493348 445352 493368
rect 445352 493348 445354 493368
rect 445298 493312 445354 493348
rect 445298 491136 445354 491192
rect 445298 487348 445354 487384
rect 445298 487328 445300 487348
rect 445300 487328 445352 487348
rect 445352 487328 445354 487348
rect 445114 441380 445170 441416
rect 445114 441360 445116 441380
rect 445116 441360 445168 441380
rect 445168 441360 445170 441380
rect 445666 509940 445668 509960
rect 445668 509940 445720 509960
rect 445720 509940 445722 509960
rect 445666 509904 445722 509940
rect 445574 509360 445630 509416
rect 445574 508816 445630 508872
rect 445666 508272 445722 508328
rect 445574 507204 445630 507240
rect 445574 507184 445576 507204
rect 445576 507184 445628 507204
rect 445628 507184 445630 507204
rect 445666 506640 445722 506696
rect 445666 506096 445722 506152
rect 445574 505552 445630 505608
rect 445666 504464 445722 504520
rect 445482 501880 445538 501936
rect 445574 500248 445630 500304
rect 445666 499704 445722 499760
rect 445574 499160 445630 499216
rect 445482 498072 445538 498128
rect 445574 497004 445630 497040
rect 445574 496984 445576 497004
rect 445576 496984 445628 497004
rect 445628 496984 445630 497004
rect 445482 488416 445538 488472
rect 445482 486240 445538 486296
rect 445482 484628 445538 484664
rect 445482 484608 445484 484628
rect 445484 484608 445536 484628
rect 445536 484608 445538 484628
rect 445574 440292 445630 440328
rect 445574 440272 445576 440292
rect 445576 440272 445628 440292
rect 445628 440272 445630 440292
rect 445574 426400 445630 426456
rect 445574 420588 445576 420608
rect 445576 420588 445628 420608
rect 445628 420588 445630 420608
rect 445574 420552 445630 420588
rect 445482 413652 445484 413672
rect 445484 413652 445536 413672
rect 445536 413652 445538 413672
rect 445482 413616 445538 413652
rect 445482 412564 445484 412584
rect 445484 412564 445536 412584
rect 445536 412564 445538 412584
rect 445482 412528 445538 412564
rect 445390 366968 445446 367024
rect 445114 363160 445170 363216
rect 445114 362072 445170 362128
rect 445114 361548 445170 361584
rect 445114 361528 445116 361548
rect 445116 361528 445168 361548
rect 445168 361528 445170 361548
rect 445114 360440 445170 360496
rect 445114 359488 445170 359544
rect 444746 358400 444802 358456
rect 444654 354592 444710 354648
rect 444378 351364 444380 351384
rect 444380 351364 444432 351384
rect 444432 351364 444434 351384
rect 444378 351328 444434 351364
rect 444378 347656 444434 347712
rect 444470 344936 444526 344992
rect 444378 343884 444380 343904
rect 444380 343884 444432 343904
rect 444432 343884 444434 343904
rect 444378 343848 444434 343884
rect 444378 297508 444380 297528
rect 444380 297508 444432 297528
rect 444432 297508 444434 297528
rect 444378 297472 444434 297508
rect 444378 296384 444434 296440
rect 443550 289448 443606 289504
rect 443182 287156 443238 287192
rect 443182 287136 443184 287156
rect 443184 287136 443236 287156
rect 443236 287136 443238 287156
rect 443090 272040 443146 272096
rect 441618 271496 441674 271552
rect 436926 265512 436982 265568
rect 434902 264968 434958 265024
rect 435178 196016 435234 196072
rect 436742 196016 436798 196072
rect 441618 226244 441620 226264
rect 441620 226244 441672 226264
rect 441672 226244 441674 226264
rect 441618 226208 441674 226244
rect 441618 225528 441674 225584
rect 441618 224868 441674 224904
rect 441618 224848 441620 224868
rect 441620 224848 441672 224868
rect 441672 224848 441674 224868
rect 441710 224440 441766 224496
rect 442078 223488 442134 223544
rect 441986 223352 442042 223408
rect 442170 221856 442226 221912
rect 442354 222400 442410 222456
rect 442262 221312 442318 221368
rect 441802 220632 441858 220688
rect 442262 211656 442318 211712
rect 442722 211656 442778 211712
rect 442170 210568 442226 210624
rect 442078 205808 442134 205864
rect 441618 204992 441674 205048
rect 441802 204584 441858 204640
rect 441710 201864 441766 201920
rect 441986 203496 442042 203552
rect 442906 205300 442908 205320
rect 442908 205300 442960 205320
rect 442960 205300 442962 205320
rect 442906 205264 442962 205300
rect 442722 203632 442778 203688
rect 442354 203088 442410 203144
rect 442906 202000 442962 202056
rect 441618 135924 441674 135960
rect 441618 135904 441620 135924
rect 441620 135904 441672 135924
rect 441672 135904 441674 135924
rect 441618 124908 441674 124944
rect 441618 124888 441620 124908
rect 441620 124888 441672 124908
rect 441672 124888 441674 124908
rect 441802 153992 441858 154048
rect 443090 219680 443146 219736
rect 443366 218592 443422 218648
rect 444286 289448 444342 289504
rect 444378 282512 444434 282568
rect 444562 340176 444618 340232
rect 444470 280064 444526 280120
rect 445022 358944 445078 359000
rect 445022 355680 445078 355736
rect 444746 284844 444802 284880
rect 444746 284824 444748 284844
rect 444748 284824 444800 284844
rect 444800 284824 444802 284844
rect 444746 281308 444802 281344
rect 444746 281288 444748 281308
rect 444748 281288 444800 281308
rect 444800 281288 444802 281308
rect 444654 277888 444710 277944
rect 444562 276664 444618 276720
rect 444562 273264 444618 273320
rect 443550 220768 443606 220824
rect 443642 219136 443698 219192
rect 443458 218048 443514 218104
rect 443274 217504 443330 217560
rect 443366 212744 443422 212800
rect 443274 212200 443330 212256
rect 443182 210024 443238 210080
rect 442998 197648 443054 197704
rect 443458 211112 443514 211168
rect 444746 274352 444802 274408
rect 444470 216008 444526 216064
rect 444378 215464 444434 215520
rect 444562 214920 444618 214976
rect 444746 223488 444802 223544
rect 444746 221856 444802 221912
rect 444746 220224 444802 220280
rect 444654 214376 444710 214432
rect 444838 213832 444894 213888
rect 444746 212200 444802 212256
rect 444286 207304 444342 207360
rect 444194 206216 444250 206272
rect 444378 205844 444380 205864
rect 444380 205844 444432 205864
rect 444432 205844 444434 205864
rect 444378 205808 444434 205844
rect 441802 151988 441804 152008
rect 441804 151988 441856 152008
rect 441856 151988 441858 152008
rect 441802 151952 441858 151988
rect 442814 158752 442870 158808
rect 442722 150320 442778 150376
rect 442262 145968 442318 146024
rect 444378 204756 444380 204776
rect 444380 204756 444432 204776
rect 444432 204756 444434 204776
rect 444378 204720 444434 204756
rect 444470 198736 444526 198792
rect 444378 147736 444434 147792
rect 443090 146512 443146 146568
rect 442998 137264 443054 137320
rect 443090 134952 443146 135008
rect 442906 129784 442962 129840
rect 441894 127472 441950 127528
rect 441802 126384 441858 126440
rect 442078 125704 442134 125760
rect 444194 132096 444250 132152
rect 444746 207848 444802 207904
rect 444838 201320 444894 201376
rect 444838 200368 444894 200424
rect 445574 364284 445576 364304
rect 445576 364284 445628 364304
rect 445628 364284 445630 364304
rect 445574 364248 445630 364284
rect 445390 360032 445446 360088
rect 445298 359488 445354 359544
rect 445206 358400 445262 358456
rect 445298 357312 445354 357368
rect 445114 353504 445170 353560
rect 445114 346604 445116 346624
rect 445116 346604 445168 346624
rect 445168 346604 445170 346624
rect 445114 346568 445170 346604
rect 445114 342252 445116 342272
rect 445116 342252 445168 342272
rect 445168 342252 445170 342272
rect 445114 342216 445170 342252
rect 445850 581984 445906 582040
rect 445758 497528 445814 497584
rect 445942 572736 445998 572792
rect 445850 495896 445906 495952
rect 445942 427488 445998 427544
rect 445666 357856 445722 357912
rect 445482 357176 445538 357232
rect 445574 356768 445630 356824
rect 445574 354068 445630 354104
rect 445574 354048 445576 354068
rect 445576 354048 445628 354068
rect 445628 354048 445630 354068
rect 445574 352960 445630 353016
rect 445574 352452 445576 352472
rect 445576 352452 445628 352472
rect 445628 352452 445630 352472
rect 445574 352416 445630 352452
rect 445574 351908 445576 351928
rect 445576 351908 445628 351928
rect 445628 351908 445630 351928
rect 445574 351872 445630 351908
rect 445482 350260 445538 350296
rect 445482 350240 445484 350260
rect 445484 350240 445536 350260
rect 445536 350240 445538 350260
rect 445482 345480 445538 345536
rect 445482 340604 445538 340640
rect 445482 340584 445484 340604
rect 445484 340584 445536 340604
rect 445536 340584 445538 340604
rect 445942 349288 445998 349344
rect 445850 347112 445906 347168
rect 445758 346024 445814 346080
rect 445390 295196 445392 295216
rect 445392 295196 445444 295216
rect 445444 295196 445446 295216
rect 445390 295160 445446 295196
rect 445482 294072 445538 294128
rect 445482 290536 445538 290592
rect 445482 280200 445538 280256
rect 445298 280064 445354 280120
rect 445298 278976 445354 279032
rect 445114 213288 445170 213344
rect 445114 212356 445170 212392
rect 445114 212336 445116 212356
rect 445116 212336 445168 212356
rect 445168 212336 445170 212356
rect 445114 209480 445170 209536
rect 445114 208392 445170 208448
rect 444930 198736 444986 198792
rect 444838 144200 444894 144256
rect 444654 140800 444710 140856
rect 444470 129784 444526 129840
rect 443366 128696 443422 128752
rect 444838 128016 444894 128072
rect 445114 206760 445170 206816
rect 445390 275576 445446 275632
rect 445206 201320 445262 201376
rect 445482 269764 445484 269784
rect 445484 269764 445536 269784
rect 445536 269764 445538 269784
rect 445482 269728 445538 269764
rect 445482 268640 445538 268696
rect 445298 201184 445354 201240
rect 445942 288224 445998 288280
rect 445850 283600 445906 283656
rect 446494 291760 446550 291816
rect 445666 222944 445722 223000
rect 445574 222400 445630 222456
rect 445574 221312 445630 221368
rect 445666 220768 445722 220824
rect 445574 219680 445630 219736
rect 445942 216960 445998 217016
rect 445850 216416 445906 216472
rect 445666 208936 445722 208992
rect 445666 207848 445722 207904
rect 445574 204176 445630 204232
rect 445206 198872 445262 198928
rect 445482 199824 445538 199880
rect 445298 198192 445354 198248
rect 445298 197648 445354 197704
rect 445022 169632 445078 169688
rect 445666 202544 445722 202600
rect 445666 201492 445668 201512
rect 445668 201492 445720 201512
rect 445720 201492 445722 201512
rect 445666 201456 445722 201492
rect 445666 197104 445722 197160
rect 445390 196560 445446 196616
rect 445850 196152 445906 196208
rect 446862 206760 446918 206816
rect 467102 354592 467158 354648
rect 449346 267688 449402 267744
rect 513378 585384 513434 585440
rect 513562 585404 513618 585440
rect 513562 585384 513564 585404
rect 513564 585384 513616 585404
rect 513616 585384 513618 585404
rect 516138 584568 516194 584624
rect 513378 583888 513434 583944
rect 513562 583888 513618 583944
rect 513378 580488 513434 580544
rect 513286 580080 513342 580136
rect 513746 582800 513802 582856
rect 513654 581712 513710 581768
rect 514850 582936 514906 582992
rect 513930 582256 513986 582312
rect 513838 580624 513894 580680
rect 513470 579536 513526 579592
rect 513470 577768 513526 577824
rect 513654 574096 513710 574152
rect 513378 556416 513434 556472
rect 513746 573552 513802 573608
rect 513930 573008 513986 573064
rect 513838 571376 513894 571432
rect 513930 556008 513986 556064
rect 513746 512660 513748 512680
rect 513748 512660 513800 512680
rect 513800 512660 513802 512680
rect 513746 512624 513802 512660
rect 513470 488688 513526 488744
rect 513378 487464 513434 487520
rect 513746 485152 513802 485208
rect 516322 578584 516378 578640
rect 516230 576952 516286 577008
rect 516690 577496 516746 577552
rect 516414 575456 516470 575512
rect 516506 572192 516562 572248
rect 516322 571104 516378 571160
rect 516230 569472 516286 569528
rect 516138 568948 516194 568984
rect 516138 568928 516140 568948
rect 516140 568928 516192 568948
rect 516192 568928 516194 568948
rect 516414 570560 516470 570616
rect 516230 567840 516286 567896
rect 516138 567316 516194 567352
rect 516138 567296 516140 567316
rect 516140 567296 516192 567316
rect 516192 567296 516194 567316
rect 516598 570016 516654 570072
rect 516506 566752 516562 566808
rect 516414 566208 516470 566264
rect 516506 565256 516562 565312
rect 516414 564712 516470 564768
rect 516322 564168 516378 564224
rect 516322 563624 516378 563680
rect 516322 563100 516378 563136
rect 516322 563080 516324 563100
rect 516324 563080 516376 563100
rect 516376 563080 516378 563100
rect 516322 562556 516378 562592
rect 516322 562536 516324 562556
rect 516324 562536 516376 562556
rect 516376 562536 516378 562556
rect 516322 562012 516378 562048
rect 516322 561992 516324 562012
rect 516324 561992 516376 562012
rect 516376 561992 516378 562012
rect 516322 561468 516378 561504
rect 516322 561448 516324 561468
rect 516324 561448 516376 561468
rect 516376 561448 516378 561468
rect 516322 559272 516378 559328
rect 516322 557676 516324 557696
rect 516324 557676 516376 557696
rect 516376 557676 516378 557696
rect 516322 557640 516378 557676
rect 516230 557096 516286 557152
rect 516138 556552 516194 556608
rect 516506 559816 516562 559872
rect 516506 558728 516562 558784
rect 516874 576408 516930 576464
rect 516782 573280 516838 573336
rect 516966 576000 517022 576056
rect 517426 574912 517482 574968
rect 517426 560904 517482 560960
rect 517242 560360 517298 560416
rect 517058 558184 517114 558240
rect 516138 512352 516194 512408
rect 516138 510040 516194 510096
rect 516138 508836 516194 508872
rect 516138 508816 516140 508836
rect 516140 508816 516192 508836
rect 516192 508816 516194 508836
rect 516138 506504 516194 506560
rect 516138 504192 516194 504248
rect 516414 507728 516470 507784
rect 516322 503104 516378 503160
rect 516138 500812 516194 500848
rect 516138 500792 516140 500812
rect 516140 500792 516192 500812
rect 516192 500792 516194 500812
rect 516138 499568 516194 499624
rect 516138 498500 516194 498536
rect 516138 498480 516140 498500
rect 516140 498480 516192 498500
rect 516192 498480 516194 498500
rect 516138 497256 516194 497312
rect 516230 496168 516286 496224
rect 516322 493856 516378 493912
rect 516230 492632 516286 492688
rect 516138 491544 516194 491600
rect 516138 490320 516194 490376
rect 516138 486920 516194 486976
rect 516138 485732 516140 485752
rect 516140 485732 516192 485752
rect 516192 485732 516194 485752
rect 516138 485696 516194 485732
rect 516690 489232 516746 489288
rect 517150 513440 517206 513496
rect 516966 505436 517022 505472
rect 516966 505416 516968 505436
rect 516968 505416 517020 505436
rect 517020 505416 517022 505436
rect 516874 501880 516930 501936
rect 516874 494944 516930 495000
rect 516138 440544 516194 440600
rect 513746 440292 513802 440328
rect 513746 440272 513748 440292
rect 513748 440272 513800 440292
rect 513800 440272 513802 440292
rect 516138 438932 516194 438968
rect 516138 438912 516140 438932
rect 516140 438912 516192 438932
rect 516192 438912 516194 438932
rect 516230 438368 516286 438424
rect 516138 437824 516194 437880
rect 516230 437280 516286 437336
rect 516138 436192 516194 436248
rect 516230 435648 516286 435704
rect 516138 435104 516194 435160
rect 516230 434016 516286 434072
rect 516138 433492 516194 433528
rect 516138 433472 516140 433492
rect 516140 433472 516192 433492
rect 516192 433472 516194 433492
rect 513470 432248 513526 432304
rect 516230 431976 516286 432032
rect 513378 430616 513434 430672
rect 516230 431432 516286 431488
rect 516506 436736 516562 436792
rect 516506 434560 516562 434616
rect 516506 432928 516562 432984
rect 516414 430888 516470 430944
rect 516414 429800 516470 429856
rect 516506 429256 516562 429312
rect 516414 428712 516470 428768
rect 516138 426536 516194 426592
rect 516322 425992 516378 426048
rect 516138 424904 516194 424960
rect 516138 424396 516140 424416
rect 516140 424396 516192 424416
rect 516192 424396 516194 424416
rect 516138 424360 516194 424396
rect 516230 423816 516286 423872
rect 516138 423272 516194 423328
rect 516322 422728 516378 422784
rect 517702 568384 517758 568440
rect 517610 565800 517666 565856
rect 517702 511128 517758 511184
rect 517426 494944 517482 495000
rect 517242 493856 517298 493912
rect 517242 488008 517298 488064
rect 516782 432384 516838 432440
rect 516874 431976 516930 432032
rect 516782 428168 516838 428224
rect 516690 427080 516746 427136
rect 517058 441632 517114 441688
rect 516966 427624 517022 427680
rect 516322 422184 516378 422240
rect 516322 421776 516378 421832
rect 516322 421232 516378 421288
rect 516322 420688 516378 420744
rect 516322 418532 516378 418568
rect 516322 418512 516324 418532
rect 516324 418512 516376 418532
rect 516376 418512 516378 418532
rect 516322 417968 516378 418024
rect 516322 415812 516378 415848
rect 516322 415792 516324 415812
rect 516324 415792 516376 415812
rect 516376 415792 516378 415812
rect 516322 414724 516378 414760
rect 516322 414704 516324 414724
rect 516324 414704 516376 414724
rect 516376 414704 516378 414724
rect 516322 414160 516378 414216
rect 516322 413072 516378 413128
rect 516322 412548 516378 412584
rect 516322 412528 516324 412548
rect 516324 412528 516376 412548
rect 516376 412528 516378 412548
rect 516506 419056 516562 419112
rect 516598 416880 516654 416936
rect 516506 416336 516562 416392
rect 516506 415248 516562 415304
rect 516782 425448 516838 425504
rect 516782 420180 516784 420200
rect 516784 420180 516836 420200
rect 516836 420180 516838 420200
rect 516782 420144 516838 420180
rect 516782 419600 516838 419656
rect 516782 413616 516838 413672
rect 445114 143112 445170 143168
rect 445298 148824 445354 148880
rect 445206 141888 445262 141944
rect 445666 152360 445722 152416
rect 445574 139576 445630 139632
rect 445298 137264 445354 137320
rect 445666 133864 445722 133920
rect 445114 132640 445170 132696
rect 445114 132096 445170 132152
rect 445942 156440 445998 156496
rect 445942 156032 445998 156088
rect 445942 151136 445998 151192
rect 445850 138488 445906 138544
rect 483662 153856 483718 153912
rect 513378 411576 513434 411632
rect 516138 369416 516194 369472
rect 513746 369164 513802 369200
rect 513746 369144 513748 369164
rect 513748 369144 513800 369164
rect 513800 369144 513802 369164
rect 516138 368364 516140 368384
rect 516140 368364 516192 368384
rect 516192 368364 516194 368384
rect 516138 368328 516194 368364
rect 513654 367940 513710 367976
rect 513654 367920 513656 367940
rect 513656 367920 513708 367940
rect 513708 367920 513710 367940
rect 513746 367648 513802 367704
rect 516138 367104 516194 367160
rect 516414 366016 516470 366072
rect 516230 364792 516286 364848
rect 516138 363704 516194 363760
rect 516138 362480 516194 362536
rect 516782 361392 516838 361448
rect 516138 360168 516194 360224
rect 516138 359116 516140 359136
rect 516140 359116 516192 359136
rect 516192 359116 516194 359136
rect 516138 359080 516194 359116
rect 516138 357892 516140 357912
rect 516140 357892 516192 357912
rect 516192 357892 516194 357912
rect 516138 357856 516194 357892
rect 516414 356768 516470 356824
rect 516138 355580 516140 355600
rect 516140 355580 516192 355600
rect 516192 355580 516194 355600
rect 516138 355544 516194 355580
rect 516138 354492 516140 354512
rect 516140 354492 516192 354512
rect 516192 354492 516194 354512
rect 516138 354456 516194 354492
rect 516138 350920 516194 350976
rect 516138 348608 516194 348664
rect 516138 347520 516194 347576
rect 516138 346316 516194 346352
rect 516138 346296 516140 346316
rect 516140 346296 516192 346316
rect 516192 346296 516194 346316
rect 516230 345208 516286 345264
rect 513378 340856 513434 340912
rect 516138 343984 516194 344040
rect 514758 342896 514814 342952
rect 516138 341708 516140 341728
rect 516140 341708 516192 341728
rect 516192 341708 516194 341728
rect 516138 341672 516194 341708
rect 516598 349852 516654 349888
rect 516598 349832 516600 349852
rect 516600 349832 516652 349852
rect 516652 349832 516654 349852
rect 513378 297472 513434 297528
rect 513378 296792 513434 296848
rect 513378 296384 513434 296440
rect 513562 296248 513618 296304
rect 513470 295840 513526 295896
rect 513378 286184 513434 286240
rect 513378 268368 513434 268424
rect 513654 287816 513710 287872
rect 513562 286728 513618 286784
rect 513930 288224 513986 288280
rect 513838 286728 513894 286784
rect 517334 441088 517390 441144
rect 517242 440000 517298 440056
rect 513746 225020 513748 225040
rect 513748 225020 513800 225040
rect 513800 225020 513802 225040
rect 513746 224984 513802 225020
rect 513746 223916 513802 223952
rect 513746 223896 513748 223916
rect 513748 223896 513800 223916
rect 513800 223896 513802 223916
rect 513378 221856 513434 221912
rect 514666 201220 514668 201240
rect 514668 201220 514720 201240
rect 514720 201220 514722 201240
rect 514666 201184 514722 201220
rect 513562 200776 513618 200832
rect 513378 199416 513434 199472
rect 514114 199996 514116 200016
rect 514116 199996 514168 200016
rect 514168 199996 514170 200016
rect 514114 199960 514170 199996
rect 514206 198872 514262 198928
rect 514114 197648 514170 197704
rect 516138 295024 516194 295080
rect 516230 294480 516286 294536
rect 516322 293936 516378 293992
rect 516230 293800 516286 293856
rect 516138 293392 516194 293448
rect 516230 292848 516286 292904
rect 516138 292304 516194 292360
rect 516322 291760 516378 291816
rect 516230 291216 516286 291272
rect 516230 290672 516286 290728
rect 516322 290128 516378 290184
rect 516138 289620 516140 289640
rect 516140 289620 516192 289640
rect 516192 289620 516194 289640
rect 516138 289584 516194 289620
rect 516230 289040 516286 289096
rect 516322 288496 516378 288552
rect 516966 297744 517022 297800
rect 516414 285368 516470 285424
rect 516782 284824 516838 284880
rect 516506 284280 516562 284336
rect 516414 283736 516470 283792
rect 516322 282648 516378 282704
rect 516138 281580 516194 281616
rect 516138 281560 516140 281580
rect 516140 281560 516192 281580
rect 516192 281560 516194 281580
rect 516230 281016 516286 281072
rect 516138 280492 516194 280528
rect 516138 280472 516140 280492
rect 516140 280472 516192 280492
rect 516192 280472 516194 280492
rect 516230 279928 516286 279984
rect 516138 279384 516194 279440
rect 516138 276820 516194 276856
rect 516138 276800 516140 276820
rect 516140 276800 516192 276820
rect 516192 276800 516194 276820
rect 516138 275204 516140 275224
rect 516140 275204 516192 275224
rect 516192 275204 516194 275224
rect 516138 275168 516194 275204
rect 516138 274660 516140 274680
rect 516140 274660 516192 274680
rect 516192 274660 516194 274680
rect 516138 274624 516194 274660
rect 516138 272992 516194 273048
rect 516138 271924 516194 271960
rect 516138 271904 516140 271924
rect 516140 271904 516192 271924
rect 516192 271904 516194 271924
rect 516138 271360 516194 271416
rect 516138 269728 516194 269784
rect 516138 269184 516194 269240
rect 516138 268660 516194 268696
rect 516138 268640 516140 268660
rect 516140 268640 516192 268660
rect 516192 268640 516194 268660
rect 516414 278296 516470 278352
rect 516322 277344 516378 277400
rect 516322 275712 516378 275768
rect 516322 272484 516324 272504
rect 516324 272484 516376 272504
rect 516376 272484 516378 272504
rect 516322 272448 516378 272484
rect 516322 270816 516378 270872
rect 516322 270272 516378 270328
rect 516598 283192 516654 283248
rect 516690 277908 516746 277944
rect 516690 277888 516692 277908
rect 516692 277888 516744 277908
rect 516744 277888 516746 277908
rect 516690 276292 516692 276312
rect 516692 276292 516744 276312
rect 516744 276292 516746 276312
rect 516690 276256 516746 276292
rect 516690 274100 516746 274136
rect 516690 274080 516692 274100
rect 516692 274080 516744 274100
rect 516744 274080 516746 274100
rect 517058 296656 517114 296712
rect 516138 225392 516194 225448
rect 516138 224304 516194 224360
rect 516138 221992 516194 222048
rect 516138 220788 516194 220824
rect 516138 220768 516140 220788
rect 516140 220768 516192 220788
rect 516192 220768 516194 220788
rect 516138 219680 516194 219736
rect 516138 218456 516194 218512
rect 516414 217368 516470 217424
rect 516138 216144 516194 216200
rect 516598 223080 516654 223136
rect 516506 215056 516562 215112
rect 516230 213868 516232 213888
rect 516232 213868 516284 213888
rect 516284 213868 516286 213888
rect 516230 213832 516286 213868
rect 516138 212744 516194 212800
rect 516138 211520 516194 211576
rect 516138 209208 516194 209264
rect 516138 206916 516194 206952
rect 516138 206896 516140 206916
rect 516140 206896 516192 206916
rect 516192 206896 516194 206916
rect 516138 205844 516140 205864
rect 516140 205844 516192 205864
rect 516192 205844 516194 205864
rect 516138 205808 516194 205844
rect 516138 204584 516194 204640
rect 516138 203496 516194 203552
rect 516138 202272 516194 202328
rect 516414 210432 516470 210488
rect 513930 156032 513986 156088
rect 513562 153856 513618 153912
rect 513378 152904 513434 152960
rect 513378 149640 513434 149696
rect 513286 148960 513342 149016
rect 513562 151680 513618 151736
rect 513470 148552 513526 148608
rect 513286 142704 513342 142760
rect 513378 134000 513434 134056
rect 513654 151272 513710 151328
rect 513838 152360 513894 152416
rect 513746 150184 513802 150240
rect 513470 132368 513526 132424
rect 513654 133592 513710 133648
rect 513930 137264 513986 137320
rect 513838 136584 513894 136640
rect 513746 133048 513802 133104
rect 513562 131416 513618 131472
rect 513286 129104 513342 129160
rect 513470 128560 513526 128616
rect 513378 125296 513434 125352
rect 513378 124888 513434 124944
rect 513838 128016 513894 128072
rect 513746 127472 513802 127528
rect 513654 125840 513710 125896
rect 513562 125296 513618 125352
rect 513286 124344 513342 124400
rect 513930 127064 513986 127120
rect 514390 151952 514446 152008
rect 514390 151816 514446 151872
rect 514206 151408 514262 151464
rect 514114 151272 514170 151328
rect 514298 150728 514354 150784
rect 514298 146104 514354 146160
rect 514298 141344 514354 141400
rect 514206 135360 514262 135416
rect 515218 141888 515274 141944
rect 515126 140800 515182 140856
rect 515034 140256 515090 140312
rect 515310 139712 515366 139768
rect 516138 152632 516194 152688
rect 516230 152088 516286 152144
rect 516322 147736 516378 147792
rect 516230 147192 516286 147248
rect 516138 145560 516194 145616
rect 516414 145016 516470 145072
rect 515586 142976 515642 143032
rect 515494 139168 515550 139224
rect 516690 146648 516746 146704
rect 516598 144472 516654 144528
rect 517426 417424 517482 417480
rect 517610 484608 517666 484664
rect 517426 352144 517482 352200
rect 517610 412120 517666 412176
rect 517610 353232 517666 353288
rect 517334 297200 517390 297256
rect 517150 282104 517206 282160
rect 517426 273536 517482 273592
rect 517794 278840 517850 278896
rect 517426 208120 517482 208176
rect 517426 196560 517482 196616
rect 516874 153720 516930 153776
rect 516782 144064 516838 144120
rect 516506 143520 516562 143576
rect 516506 138624 516562 138680
rect 516230 138080 516286 138136
rect 516138 137536 516194 137592
rect 514942 135904 514998 135960
rect 514850 134816 514906 134872
rect 514758 134272 514814 134328
rect 514114 131688 514170 131744
rect 516138 130600 516194 130656
rect 514114 126384 514170 126440
rect 516230 130056 516286 130112
rect 517426 124208 517482 124264
rect 517610 153176 517666 153232
rect 450542 97416 450598 97472
rect 447782 97280 447838 97336
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580262 577632 580318 577688
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 325216 579674 325272
rect 580170 312024 580226 312080
rect 580354 564304 580410 564360
rect 582378 511264 582434 511320
rect 580446 431568 580502 431624
rect 580538 418240 580594 418296
rect 580630 365064 580686 365120
rect 580722 351872 580778 351928
rect 582470 484608 582526 484664
rect 580170 298696 580226 298752
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 272176 580502 272232
rect 580354 258848 580410 258904
rect 580262 232328 580318 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 532698 95920 532754 95976
rect 547142 95784 547198 95840
rect 580262 97144 580318 97200
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 582470 46280 582526 46336
rect 582378 6568 582434 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 371233 585714 371299 585717
rect 369932 585712 371299 585714
rect 369932 585656 371238 585712
rect 371294 585656 371299 585712
rect 369932 585654 371299 585656
rect 371233 585651 371299 585654
rect 513422 585445 513482 585684
rect 445661 585442 445727 585445
rect 441876 585440 445727 585442
rect 441876 585384 445666 585440
rect 445722 585384 445727 585440
rect 441876 585382 445727 585384
rect 445661 585379 445727 585382
rect 513373 585440 513482 585445
rect 513373 585384 513378 585440
rect 513434 585384 513482 585440
rect 513373 585382 513482 585384
rect 513557 585442 513623 585445
rect 513557 585440 513666 585442
rect 513557 585384 513562 585440
rect 513618 585384 513666 585440
rect 513373 585379 513439 585382
rect 513557 585379 513666 585384
rect 371693 585170 371759 585173
rect 369932 585168 371759 585170
rect 369932 585112 371698 585168
rect 371754 585112 371759 585168
rect 513606 585140 513666 585379
rect 369932 585110 371759 585112
rect 371693 585107 371759 585110
rect 371417 584626 371483 584629
rect 516133 584626 516199 584629
rect 369932 584624 371483 584626
rect 369932 584568 371422 584624
rect 371478 584568 371483 584624
rect 369932 584566 371483 584568
rect 513820 584624 516199 584626
rect 513820 584568 516138 584624
rect 516194 584568 516199 584624
rect 513820 584566 516199 584568
rect 371417 584563 371483 584566
rect 516133 584563 516199 584566
rect 444741 584354 444807 584357
rect 441876 584352 444807 584354
rect 441876 584296 444746 584352
rect 444802 584296 444807 584352
rect 441876 584294 444807 584296
rect 444741 584291 444807 584294
rect 371182 584082 371188 584084
rect 369932 584022 371188 584082
rect 371182 584020 371188 584022
rect 371252 584020 371258 584084
rect 513422 583949 513482 584052
rect 513373 583944 513482 583949
rect 513373 583888 513378 583944
rect 513434 583888 513482 583944
rect 513373 583886 513482 583888
rect 513557 583946 513623 583949
rect 513557 583944 513666 583946
rect 513557 583888 513562 583944
rect 513618 583888 513666 583944
rect 513373 583883 513439 583886
rect 513557 583883 513666 583888
rect 371366 583538 371372 583540
rect 369932 583478 371372 583538
rect 371366 583476 371372 583478
rect 371436 583476 371442 583540
rect 513606 583508 513666 583883
rect 442993 583130 443059 583133
rect 441876 583128 443059 583130
rect 441876 583072 442998 583128
rect 443054 583072 443059 583128
rect 441876 583070 443059 583072
rect 442993 583067 443059 583070
rect 371550 582994 371556 582996
rect 369932 582934 371556 582994
rect 371550 582932 371556 582934
rect 371620 582932 371626 582996
rect 514845 582994 514911 582997
rect 513820 582992 514911 582994
rect 513820 582936 514850 582992
rect 514906 582936 514911 582992
rect 513820 582934 514911 582936
rect 514845 582931 514911 582934
rect 513741 582858 513807 582861
rect 513741 582856 513850 582858
rect 513741 582800 513746 582856
rect 513802 582800 513850 582856
rect 513741 582795 513850 582800
rect 371785 582450 371851 582453
rect 372153 582450 372219 582453
rect 369932 582448 372219 582450
rect 369932 582392 371790 582448
rect 371846 582392 372158 582448
rect 372214 582392 372219 582448
rect 513790 582420 513850 582795
rect 369932 582390 372219 582392
rect 371785 582387 371851 582390
rect 372153 582387 372219 582390
rect 513925 582314 513991 582317
rect 513790 582312 513991 582314
rect 513790 582256 513930 582312
rect 513986 582256 513991 582312
rect 513790 582254 513991 582256
rect 445845 582042 445911 582045
rect 441876 582040 445911 582042
rect 441876 581984 445850 582040
rect 445906 581984 445911 582040
rect 441876 581982 445911 581984
rect 445845 581979 445911 581982
rect 371325 581906 371391 581909
rect 369932 581904 371391 581906
rect 369932 581848 371330 581904
rect 371386 581848 371391 581904
rect 513790 581876 513850 582254
rect 513925 582251 513991 582254
rect 369932 581846 371391 581848
rect 371325 581843 371391 581846
rect 513649 581770 513715 581773
rect 513606 581768 513715 581770
rect 513606 581712 513654 581768
rect 513710 581712 513715 581768
rect 513606 581707 513715 581712
rect 371601 581362 371667 581365
rect 369932 581360 371667 581362
rect 369932 581304 371606 581360
rect 371662 581304 371667 581360
rect 513606 581332 513666 581707
rect 369932 581302 371667 581304
rect 371601 581299 371667 581302
rect 371693 580818 371759 580821
rect 443085 580818 443151 580821
rect 369932 580816 371759 580818
rect 369932 580760 371698 580816
rect 371754 580760 371759 580816
rect 369932 580758 371759 580760
rect 441876 580816 443151 580818
rect 441876 580760 443090 580816
rect 443146 580760 443151 580816
rect 441876 580758 443151 580760
rect 371693 580755 371759 580758
rect 443085 580755 443151 580758
rect 513422 580549 513482 580788
rect 513833 580682 513899 580685
rect 513373 580544 513482 580549
rect 513373 580488 513378 580544
rect 513434 580488 513482 580544
rect 513373 580486 513482 580488
rect 513790 580680 513899 580682
rect 513790 580624 513838 580680
rect 513894 580624 513899 580680
rect 513790 580619 513899 580624
rect 513373 580483 513439 580486
rect 371509 580274 371575 580277
rect 369932 580272 371575 580274
rect 369932 580216 371514 580272
rect 371570 580216 371575 580272
rect 513790 580244 513850 580619
rect 369932 580214 371575 580216
rect 371509 580211 371575 580214
rect 513281 580138 513347 580141
rect 513281 580136 513482 580138
rect -960 580002 480 580092
rect 513281 580080 513286 580136
rect 513342 580080 513482 580136
rect 513281 580078 513482 580080
rect 513281 580075 513347 580078
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 371601 579730 371667 579733
rect 444741 579730 444807 579733
rect 369932 579728 371667 579730
rect 369932 579672 371606 579728
rect 371662 579672 371667 579728
rect 369932 579670 371667 579672
rect 441876 579728 444807 579730
rect 441876 579672 444746 579728
rect 444802 579672 444807 579728
rect 513422 579700 513482 580078
rect 441876 579670 444807 579672
rect 371601 579667 371667 579670
rect 444741 579667 444807 579670
rect 513465 579594 513531 579597
rect 513422 579592 513531 579594
rect 513422 579536 513470 579592
rect 513526 579536 513531 579592
rect 513422 579531 513531 579536
rect 371693 579186 371759 579189
rect 369932 579184 371759 579186
rect 369932 579128 371698 579184
rect 371754 579128 371759 579184
rect 513422 579156 513482 579531
rect 369932 579126 371759 579128
rect 371693 579123 371759 579126
rect 371325 578642 371391 578645
rect 516317 578642 516383 578645
rect 369932 578640 371391 578642
rect 369932 578584 371330 578640
rect 371386 578584 371391 578640
rect 369932 578582 371391 578584
rect 513820 578640 516383 578642
rect 513820 578584 516322 578640
rect 516378 578584 516383 578640
rect 513820 578582 516383 578584
rect 371325 578579 371391 578582
rect 516317 578579 516383 578582
rect 444925 578506 444991 578509
rect 441876 578504 444991 578506
rect 441876 578448 444930 578504
rect 444986 578448 444991 578504
rect 441876 578446 444991 578448
rect 444925 578443 444991 578446
rect 371693 578098 371759 578101
rect 369932 578096 371759 578098
rect 369932 578040 371698 578096
rect 371754 578040 371759 578096
rect 369932 578038 371759 578040
rect 371693 578035 371759 578038
rect 513422 577829 513482 578068
rect 513422 577824 513531 577829
rect 513422 577768 513470 577824
rect 513526 577768 513531 577824
rect 513422 577766 513531 577768
rect 513465 577763 513531 577766
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 371417 577554 371483 577557
rect 516685 577554 516751 577557
rect 369932 577552 371483 577554
rect 369932 577496 371422 577552
rect 371478 577496 371483 577552
rect 369932 577494 371483 577496
rect 513820 577552 516751 577554
rect 513820 577496 516690 577552
rect 516746 577496 516751 577552
rect 583520 577540 584960 577630
rect 513820 577494 516751 577496
rect 371417 577491 371483 577494
rect 516685 577491 516751 577494
rect 441662 577149 441722 577388
rect 441613 577144 441722 577149
rect 441613 577088 441618 577144
rect 441674 577088 441722 577144
rect 441613 577086 441722 577088
rect 441613 577083 441679 577086
rect 371601 577010 371667 577013
rect 516225 577010 516291 577013
rect 369932 577008 371667 577010
rect 369932 576952 371606 577008
rect 371662 576952 371667 577008
rect 369932 576950 371667 576952
rect 513820 577008 516291 577010
rect 513820 576952 516230 577008
rect 516286 576952 516291 577008
rect 513820 576950 516291 576952
rect 371601 576947 371667 576950
rect 516225 576947 516291 576950
rect 371693 576466 371759 576469
rect 516869 576466 516935 576469
rect 369932 576464 371759 576466
rect 369932 576408 371698 576464
rect 371754 576408 371759 576464
rect 369932 576406 371759 576408
rect 513820 576464 516935 576466
rect 513820 576408 516874 576464
rect 516930 576408 516935 576464
rect 513820 576406 516935 576408
rect 371693 576403 371759 576406
rect 516869 576403 516935 576406
rect 444741 576194 444807 576197
rect 441876 576192 444807 576194
rect 441876 576136 444746 576192
rect 444802 576136 444807 576192
rect 441876 576134 444807 576136
rect 444741 576131 444807 576134
rect 371877 576058 371943 576061
rect 516961 576058 517027 576061
rect 369932 576056 371943 576058
rect 369932 576000 371882 576056
rect 371938 576000 371943 576056
rect 369932 575998 371943 576000
rect 513820 576056 517027 576058
rect 513820 576000 516966 576056
rect 517022 576000 517027 576056
rect 513820 575998 517027 576000
rect 371877 575995 371943 575998
rect 516961 575995 517027 575998
rect 371601 575514 371667 575517
rect 516409 575514 516475 575517
rect 369932 575512 371667 575514
rect 369932 575456 371606 575512
rect 371662 575456 371667 575512
rect 369932 575454 371667 575456
rect 513820 575512 516475 575514
rect 513820 575456 516414 575512
rect 516470 575456 516475 575512
rect 513820 575454 516475 575456
rect 371601 575451 371667 575454
rect 516409 575451 516475 575454
rect 444557 575106 444623 575109
rect 441876 575104 444623 575106
rect 441876 575048 444562 575104
rect 444618 575048 444623 575104
rect 441876 575046 444623 575048
rect 444557 575043 444623 575046
rect 371785 574970 371851 574973
rect 517421 574970 517487 574973
rect 369932 574968 371851 574970
rect 369932 574912 371790 574968
rect 371846 574912 371851 574968
rect 369932 574910 371851 574912
rect 513820 574968 517487 574970
rect 513820 574912 517426 574968
rect 517482 574912 517487 574968
rect 513820 574910 517487 574912
rect 371785 574907 371851 574910
rect 517421 574907 517487 574910
rect 372429 574426 372495 574429
rect 369932 574424 372495 574426
rect 369932 574368 372434 574424
rect 372490 574368 372495 574424
rect 369932 574366 372495 574368
rect 372429 574363 372495 574366
rect 513606 574157 513666 574396
rect 513606 574152 513715 574157
rect 513606 574096 513654 574152
rect 513710 574096 513715 574152
rect 513606 574094 513715 574096
rect 513649 574091 513715 574094
rect 371969 573882 372035 573885
rect 369932 573880 372035 573882
rect 369932 573824 371974 573880
rect 372030 573824 372035 573880
rect 369932 573822 372035 573824
rect 371969 573819 372035 573822
rect 441846 573341 441906 573852
rect 513790 573613 513850 573852
rect 513741 573608 513850 573613
rect 513741 573552 513746 573608
rect 513802 573552 513850 573608
rect 513741 573550 513850 573552
rect 513741 573547 513807 573550
rect 372061 573338 372127 573341
rect 369932 573336 372127 573338
rect 369932 573280 372066 573336
rect 372122 573280 372127 573336
rect 369932 573278 372127 573280
rect 372061 573275 372127 573278
rect 441797 573336 441906 573341
rect 516777 573338 516843 573341
rect 441797 573280 441802 573336
rect 441858 573280 441906 573336
rect 441797 573278 441906 573280
rect 513820 573336 516843 573338
rect 513820 573280 516782 573336
rect 516838 573280 516843 573336
rect 513820 573278 516843 573280
rect 441797 573275 441863 573278
rect 516777 573275 516843 573278
rect 513925 573066 513991 573069
rect 513790 573064 513991 573066
rect 513790 573008 513930 573064
rect 513986 573008 513991 573064
rect 513790 573006 513991 573008
rect 372245 572794 372311 572797
rect 445937 572794 446003 572797
rect 369932 572792 372311 572794
rect 369932 572736 372250 572792
rect 372306 572736 372311 572792
rect 369932 572734 372311 572736
rect 441876 572792 446003 572794
rect 441876 572736 445942 572792
rect 445998 572736 446003 572792
rect 513790 572764 513850 573006
rect 513925 573003 513991 573006
rect 441876 572734 446003 572736
rect 372245 572731 372311 572734
rect 445937 572731 446003 572734
rect 371734 572250 371740 572252
rect 369932 572190 371740 572250
rect 371734 572188 371740 572190
rect 371804 572188 371810 572252
rect 516501 572250 516567 572253
rect 513820 572248 516567 572250
rect 513820 572192 516506 572248
rect 516562 572192 516567 572248
rect 513820 572190 516567 572192
rect 516501 572187 516567 572190
rect 371601 571706 371667 571709
rect 369932 571704 371667 571706
rect 369932 571648 371606 571704
rect 371662 571648 371667 571704
rect 369932 571646 371667 571648
rect 371601 571643 371667 571646
rect 444833 571570 444899 571573
rect 441876 571568 444899 571570
rect 441876 571512 444838 571568
rect 444894 571512 444899 571568
rect 441876 571510 444899 571512
rect 444833 571507 444899 571510
rect 513790 571437 513850 571676
rect 513790 571432 513899 571437
rect 513790 571376 513838 571432
rect 513894 571376 513899 571432
rect 513790 571374 513899 571376
rect 513833 571371 513899 571374
rect 371693 571162 371759 571165
rect 516317 571162 516383 571165
rect 369932 571160 371759 571162
rect 369932 571104 371698 571160
rect 371754 571104 371759 571160
rect 369932 571102 371759 571104
rect 513820 571160 516383 571162
rect 513820 571104 516322 571160
rect 516378 571104 516383 571160
rect 513820 571102 516383 571104
rect 371693 571099 371759 571102
rect 516317 571099 516383 571102
rect 371509 570618 371575 570621
rect 516409 570618 516475 570621
rect 369932 570616 371575 570618
rect 369932 570560 371514 570616
rect 371570 570560 371575 570616
rect 369932 570558 371575 570560
rect 513820 570616 516475 570618
rect 513820 570560 516414 570616
rect 516470 570560 516475 570616
rect 513820 570558 516475 570560
rect 371509 570555 371575 570558
rect 516409 570555 516475 570558
rect 443177 570482 443243 570485
rect 441876 570480 443243 570482
rect 441876 570424 443182 570480
rect 443238 570424 443243 570480
rect 441876 570422 443243 570424
rect 443177 570419 443243 570422
rect 371601 570074 371667 570077
rect 516593 570074 516659 570077
rect 369932 570072 371667 570074
rect 369932 570016 371606 570072
rect 371662 570016 371667 570072
rect 369932 570014 371667 570016
rect 513820 570072 516659 570074
rect 513820 570016 516598 570072
rect 516654 570016 516659 570072
rect 513820 570014 516659 570016
rect 371601 570011 371667 570014
rect 516593 570011 516659 570014
rect 516225 569530 516291 569533
rect 513820 569528 516291 569530
rect 369902 569261 369962 569500
rect 513820 569472 516230 569528
rect 516286 569472 516291 569528
rect 513820 569470 516291 569472
rect 516225 569467 516291 569470
rect 369853 569256 369962 569261
rect 444925 569258 444991 569261
rect 369853 569200 369858 569256
rect 369914 569200 369962 569256
rect 369853 569198 369962 569200
rect 441876 569256 444991 569258
rect 441876 569200 444930 569256
rect 444986 569200 444991 569256
rect 441876 569198 444991 569200
rect 369853 569195 369919 569198
rect 444925 569195 444991 569198
rect 516133 568986 516199 568989
rect 513820 568984 516199 568986
rect 369350 568717 369410 568956
rect 513820 568928 516138 568984
rect 516194 568928 516199 568984
rect 513820 568926 516199 568928
rect 516133 568923 516199 568926
rect 369301 568712 369410 568717
rect 369301 568656 369306 568712
rect 369362 568656 369410 568712
rect 369301 568654 369410 568656
rect 369301 568651 369367 568654
rect 371509 568442 371575 568445
rect 517697 568442 517763 568445
rect 369932 568440 371575 568442
rect 369932 568384 371514 568440
rect 371570 568384 371575 568440
rect 369932 568382 371575 568384
rect 513820 568440 517763 568442
rect 513820 568384 517702 568440
rect 517758 568384 517763 568440
rect 513820 568382 517763 568384
rect 371509 568379 371575 568382
rect 517697 568379 517763 568382
rect 371601 567898 371667 567901
rect 369932 567896 371667 567898
rect 369932 567840 371606 567896
rect 371662 567840 371667 567896
rect 369932 567838 371667 567840
rect 371601 567835 371667 567838
rect 441846 567629 441906 568140
rect 516225 567898 516291 567901
rect 513820 567896 516291 567898
rect 513820 567840 516230 567896
rect 516286 567840 516291 567896
rect 513820 567838 516291 567840
rect 516225 567835 516291 567838
rect 441846 567624 441955 567629
rect 441846 567568 441894 567624
rect 441950 567568 441955 567624
rect 441846 567566 441955 567568
rect 441889 567563 441955 567566
rect 516133 567354 516199 567357
rect 513820 567352 516199 567354
rect 369902 567221 369962 567324
rect 513820 567296 516138 567352
rect 516194 567296 516199 567352
rect 513820 567294 516199 567296
rect 516133 567291 516199 567294
rect 369902 567216 370011 567221
rect 369902 567160 369950 567216
rect 370006 567160 370011 567216
rect 369902 567158 370011 567160
rect 369945 567155 370011 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect 443269 566946 443335 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect 441876 566944 443335 566946
rect 441876 566888 443274 566944
rect 443330 566888 443335 566944
rect 441876 566886 443335 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 443269 566883 443335 566886
rect 516501 566810 516567 566813
rect 513820 566808 516567 566810
rect 369350 566541 369410 566780
rect 513820 566752 516506 566808
rect 516562 566752 516567 566808
rect 513820 566750 516567 566752
rect 516501 566747 516567 566750
rect 369301 566536 369410 566541
rect 369301 566480 369306 566536
rect 369362 566480 369410 566536
rect 369301 566478 369410 566480
rect 369301 566475 369367 566478
rect 371785 566266 371851 566269
rect 516409 566266 516475 566269
rect 369932 566264 371851 566266
rect 369932 566208 371790 566264
rect 371846 566208 371851 566264
rect 369932 566206 371851 566208
rect 513820 566264 516475 566266
rect 513820 566208 516414 566264
rect 516470 566208 516475 566264
rect 513820 566206 516475 566208
rect 371785 566203 371851 566206
rect 516409 566203 516475 566206
rect 371785 565858 371851 565861
rect 444465 565858 444531 565861
rect 517605 565858 517671 565861
rect 369932 565856 371851 565858
rect 369932 565800 371790 565856
rect 371846 565800 371851 565856
rect 369932 565798 371851 565800
rect 441876 565856 444531 565858
rect 441876 565800 444470 565856
rect 444526 565800 444531 565856
rect 441876 565798 444531 565800
rect 513820 565856 517671 565858
rect 513820 565800 517610 565856
rect 517666 565800 517671 565856
rect 513820 565798 517671 565800
rect 371785 565795 371851 565798
rect 444465 565795 444531 565798
rect 517605 565795 517671 565798
rect 372521 565314 372587 565317
rect 516501 565314 516567 565317
rect 369932 565312 372587 565314
rect 369932 565256 372526 565312
rect 372582 565256 372587 565312
rect 369932 565254 372587 565256
rect 513820 565312 516567 565314
rect 513820 565256 516506 565312
rect 516562 565256 516567 565312
rect 513820 565254 516567 565256
rect 372521 565251 372587 565254
rect 516501 565251 516567 565254
rect 371785 564770 371851 564773
rect 516409 564770 516475 564773
rect 369932 564768 371851 564770
rect 369932 564712 371790 564768
rect 371846 564712 371851 564768
rect 369932 564710 371851 564712
rect 513820 564768 516475 564770
rect 513820 564712 516414 564768
rect 516470 564712 516475 564768
rect 513820 564710 516475 564712
rect 371785 564707 371851 564710
rect 516409 564707 516475 564710
rect 444373 564634 444439 564637
rect 441876 564632 444439 564634
rect 441876 564576 444378 564632
rect 444434 564576 444439 564632
rect 441876 564574 444439 564576
rect 444373 564571 444439 564574
rect 580349 564362 580415 564365
rect 583520 564362 584960 564452
rect 580349 564360 584960 564362
rect 580349 564304 580354 564360
rect 580410 564304 584960 564360
rect 580349 564302 584960 564304
rect 580349 564299 580415 564302
rect 370129 564226 370195 564229
rect 516317 564226 516383 564229
rect 369932 564224 370195 564226
rect 369932 564168 370134 564224
rect 370190 564168 370195 564224
rect 369932 564166 370195 564168
rect 513820 564224 516383 564226
rect 513820 564168 516322 564224
rect 516378 564168 516383 564224
rect 583520 564212 584960 564302
rect 513820 564166 516383 564168
rect 370129 564163 370195 564166
rect 516317 564163 516383 564166
rect 372705 563682 372771 563685
rect 516317 563682 516383 563685
rect 369932 563680 372771 563682
rect 369932 563624 372710 563680
rect 372766 563624 372771 563680
rect 369932 563622 372771 563624
rect 513820 563680 516383 563682
rect 513820 563624 516322 563680
rect 516378 563624 516383 563680
rect 513820 563622 516383 563624
rect 372705 563619 372771 563622
rect 516317 563619 516383 563622
rect 445661 563546 445727 563549
rect 441876 563544 445727 563546
rect 441876 563488 445666 563544
rect 445722 563488 445727 563544
rect 441876 563486 445727 563488
rect 445661 563483 445727 563486
rect 371785 563138 371851 563141
rect 516317 563138 516383 563141
rect 369932 563136 371851 563138
rect 369932 563080 371790 563136
rect 371846 563080 371851 563136
rect 369932 563078 371851 563080
rect 513820 563136 516383 563138
rect 513820 563080 516322 563136
rect 516378 563080 516383 563136
rect 513820 563078 516383 563080
rect 371785 563075 371851 563078
rect 516317 563075 516383 563078
rect 371785 562594 371851 562597
rect 516317 562594 516383 562597
rect 369932 562592 371851 562594
rect 369932 562536 371790 562592
rect 371846 562536 371851 562592
rect 369932 562534 371851 562536
rect 513820 562592 516383 562594
rect 513820 562536 516322 562592
rect 516378 562536 516383 562592
rect 513820 562534 516383 562536
rect 371785 562531 371851 562534
rect 516317 562531 516383 562534
rect 370221 562050 370287 562053
rect 369932 562048 370287 562050
rect 369932 561992 370226 562048
rect 370282 561992 370287 562048
rect 369932 561990 370287 561992
rect 370221 561987 370287 561990
rect 441846 561778 441906 562292
rect 516317 562050 516383 562053
rect 513820 562048 516383 562050
rect 513820 561992 516322 562048
rect 516378 561992 516383 562048
rect 513820 561990 516383 561992
rect 516317 561987 516383 561990
rect 441981 561778 442047 561781
rect 441846 561776 442047 561778
rect 441846 561720 441986 561776
rect 442042 561720 442047 561776
rect 441846 561718 442047 561720
rect 441981 561715 442047 561718
rect 370313 561506 370379 561509
rect 516317 561506 516383 561509
rect 369932 561504 370379 561506
rect 369932 561448 370318 561504
rect 370374 561448 370379 561504
rect 369932 561446 370379 561448
rect 513820 561504 516383 561506
rect 513820 561448 516322 561504
rect 516378 561448 516383 561504
rect 513820 561446 516383 561448
rect 370313 561443 370379 561446
rect 516317 561443 516383 561446
rect 444373 561234 444439 561237
rect 441876 561232 444439 561234
rect 441876 561176 444378 561232
rect 444434 561176 444439 561232
rect 441876 561174 444439 561176
rect 444373 561171 444439 561174
rect 371785 560962 371851 560965
rect 517421 560962 517487 560965
rect 369932 560960 371851 560962
rect 369932 560904 371790 560960
rect 371846 560904 371851 560960
rect 369932 560902 371851 560904
rect 513820 560960 517487 560962
rect 513820 560904 517426 560960
rect 517482 560904 517487 560960
rect 513820 560902 517487 560904
rect 371785 560899 371851 560902
rect 517421 560899 517487 560902
rect 371785 560418 371851 560421
rect 517237 560418 517303 560421
rect 369932 560416 371851 560418
rect 369932 560360 371790 560416
rect 371846 560360 371851 560416
rect 369932 560358 371851 560360
rect 513820 560416 517303 560418
rect 513820 560360 517242 560416
rect 517298 560360 517303 560416
rect 513820 560358 517303 560360
rect 371785 560355 371851 560358
rect 517237 560355 517303 560358
rect 371877 559874 371943 559877
rect 369932 559872 371943 559874
rect 369932 559816 371882 559872
rect 371938 559816 371943 559872
rect 369932 559814 371943 559816
rect 371877 559811 371943 559814
rect 441662 559469 441722 559980
rect 516501 559874 516567 559877
rect 513820 559872 516567 559874
rect 513820 559816 516506 559872
rect 516562 559816 516567 559872
rect 513820 559814 516567 559816
rect 516501 559811 516567 559814
rect 441613 559464 441722 559469
rect 441613 559408 441618 559464
rect 441674 559408 441722 559464
rect 441613 559406 441722 559408
rect 441613 559403 441679 559406
rect 371785 559330 371851 559333
rect 516317 559330 516383 559333
rect 369932 559328 371851 559330
rect 369932 559272 371790 559328
rect 371846 559272 371851 559328
rect 369932 559270 371851 559272
rect 513820 559328 516383 559330
rect 513820 559272 516322 559328
rect 516378 559272 516383 559328
rect 513820 559270 516383 559272
rect 371785 559267 371851 559270
rect 516317 559267 516383 559270
rect 442073 558922 442139 558925
rect 441876 558920 442139 558922
rect 441876 558864 442078 558920
rect 442134 558864 442139 558920
rect 441876 558862 442139 558864
rect 442073 558859 442139 558862
rect 371785 558786 371851 558789
rect 516501 558786 516567 558789
rect 369932 558784 371851 558786
rect 369932 558728 371790 558784
rect 371846 558728 371851 558784
rect 369932 558726 371851 558728
rect 513820 558784 516567 558786
rect 513820 558728 516506 558784
rect 516562 558728 516567 558784
rect 513820 558726 516567 558728
rect 371785 558723 371851 558726
rect 516501 558723 516567 558726
rect 370405 558242 370471 558245
rect 517053 558242 517119 558245
rect 369932 558240 370471 558242
rect 369932 558184 370410 558240
rect 370466 558184 370471 558240
rect 369932 558182 370471 558184
rect 513820 558240 517119 558242
rect 513820 558184 517058 558240
rect 517114 558184 517119 558240
rect 513820 558182 517119 558184
rect 370405 558179 370471 558182
rect 517053 558179 517119 558182
rect 371785 557698 371851 557701
rect 444373 557698 444439 557701
rect 516317 557698 516383 557701
rect 369932 557696 371851 557698
rect 369932 557640 371790 557696
rect 371846 557640 371851 557696
rect 369932 557638 371851 557640
rect 441876 557696 444439 557698
rect 441876 557640 444378 557696
rect 444434 557640 444439 557696
rect 441876 557638 444439 557640
rect 513820 557696 516383 557698
rect 513820 557640 516322 557696
rect 516378 557640 516383 557696
rect 513820 557638 516383 557640
rect 371785 557635 371851 557638
rect 444373 557635 444439 557638
rect 516317 557635 516383 557638
rect 372797 557154 372863 557157
rect 516225 557154 516291 557157
rect 369932 557152 372863 557154
rect 369932 557096 372802 557152
rect 372858 557096 372863 557152
rect 369932 557094 372863 557096
rect 513820 557152 516291 557154
rect 513820 557096 516230 557152
rect 516286 557096 516291 557152
rect 513820 557094 516291 557096
rect 372797 557091 372863 557094
rect 516225 557091 516291 557094
rect 441705 556882 441771 556885
rect 441662 556880 441771 556882
rect 441662 556824 441710 556880
rect 441766 556824 441771 556880
rect 441662 556819 441771 556824
rect 371785 556610 371851 556613
rect 369932 556608 371851 556610
rect 369932 556552 371790 556608
rect 371846 556552 371851 556608
rect 441662 556580 441722 556819
rect 516133 556610 516199 556613
rect 513820 556608 516199 556610
rect 369932 556550 371851 556552
rect 513820 556552 516138 556608
rect 516194 556552 516199 556608
rect 513820 556550 516199 556552
rect 371785 556547 371851 556550
rect 516133 556547 516199 556550
rect 513373 556474 513439 556477
rect 513373 556472 513482 556474
rect 513373 556416 513378 556472
rect 513434 556416 513482 556472
rect 513373 556411 513482 556416
rect 370497 556202 370563 556205
rect 369932 556200 370563 556202
rect 369932 556144 370502 556200
rect 370558 556144 370563 556200
rect 513422 556172 513482 556411
rect 369932 556142 370563 556144
rect 370497 556139 370563 556142
rect 372245 556066 372311 556069
rect 513925 556066 513991 556069
rect 372245 556064 513991 556066
rect 372245 556008 372250 556064
rect 372306 556008 513930 556064
rect 513986 556008 513991 556064
rect 372245 556006 513991 556008
rect 372245 556003 372311 556006
rect 513925 556003 513991 556006
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 361614 553420 361620 553484
rect 361684 553482 361690 553484
rect 362861 553482 362927 553485
rect 361684 553480 362927 553482
rect 361684 553424 362866 553480
rect 362922 553424 362927 553480
rect 361684 553422 362927 553424
rect 361684 553420 361690 553422
rect 362861 553419 362927 553422
rect 364885 553482 364951 553485
rect 435173 553484 435239 553485
rect 436737 553484 436803 553485
rect 365294 553482 365300 553484
rect 364885 553480 365300 553482
rect 364885 553424 364890 553480
rect 364946 553424 365300 553480
rect 364885 553422 365300 553424
rect 364885 553419 364951 553422
rect 365294 553420 365300 553422
rect 365364 553420 365370 553484
rect 435173 553482 435220 553484
rect 435128 553480 435220 553482
rect 435128 553424 435178 553480
rect 435128 553422 435220 553424
rect 435173 553420 435220 553422
rect 435284 553420 435290 553484
rect 436686 553482 436692 553484
rect 436646 553422 436692 553482
rect 436756 553480 436803 553484
rect 436798 553424 436803 553480
rect 436686 553420 436692 553422
rect 436756 553420 436803 553424
rect 435173 553419 435239 553420
rect 436737 553419 436803 553420
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 444373 513770 444439 513773
rect 441876 513768 444439 513770
rect 441876 513712 444378 513768
rect 444434 513712 444439 513768
rect 441876 513710 444439 513712
rect 444373 513707 444439 513710
rect 517145 513498 517211 513501
rect 513820 513496 517211 513498
rect 369902 512957 369962 513468
rect 513820 513440 517150 513496
rect 517206 513440 517211 513496
rect 513820 513438 517211 513440
rect 517145 513435 517211 513438
rect 444833 513226 444899 513229
rect 441876 513224 444899 513226
rect 441876 513168 444838 513224
rect 444894 513168 444899 513224
rect 441876 513166 444899 513168
rect 444833 513163 444899 513166
rect 369853 512952 369962 512957
rect 369853 512896 369858 512952
rect 369914 512896 369962 512952
rect 369853 512894 369962 512896
rect 369853 512891 369919 512894
rect 444373 512682 444439 512685
rect 441876 512680 444439 512682
rect 441876 512624 444378 512680
rect 444434 512624 444439 512680
rect 441876 512622 444439 512624
rect 444373 512619 444439 512622
rect 513741 512682 513807 512685
rect 513741 512680 513850 512682
rect 513741 512624 513746 512680
rect 513802 512624 513850 512680
rect 513741 512619 513850 512624
rect 513790 512410 513850 512619
rect 516133 512410 516199 512413
rect 513790 512408 516199 512410
rect 513790 512380 516138 512408
rect 369350 511869 369410 512380
rect 513820 512352 516138 512380
rect 516194 512352 516199 512408
rect 513820 512350 516199 512352
rect 516133 512347 516199 512350
rect 444557 512138 444623 512141
rect 441876 512136 444623 512138
rect 441876 512080 444562 512136
rect 444618 512080 444623 512136
rect 441876 512078 444623 512080
rect 444557 512075 444623 512078
rect 369350 511864 369459 511869
rect 369350 511808 369398 511864
rect 369454 511808 369459 511864
rect 369350 511806 369459 511808
rect 369393 511803 369459 511806
rect 444598 511594 444604 511596
rect 441876 511534 444604 511594
rect 444598 511532 444604 511534
rect 444668 511594 444674 511596
rect 445661 511594 445727 511597
rect 444668 511592 445727 511594
rect 444668 511536 445666 511592
rect 445722 511536 445727 511592
rect 444668 511534 445727 511536
rect 444668 511532 444674 511534
rect 445661 511531 445727 511534
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 370957 511186 371023 511189
rect 517697 511186 517763 511189
rect 369932 511184 371023 511186
rect 369932 511128 370962 511184
rect 371018 511128 371023 511184
rect 369932 511126 371023 511128
rect 513820 511184 517763 511186
rect 513820 511128 517702 511184
rect 517758 511128 517763 511184
rect 583520 511172 584960 511262
rect 513820 511126 517763 511128
rect 370957 511123 371023 511126
rect 517697 511123 517763 511126
rect 445385 511050 445451 511053
rect 441876 511048 445451 511050
rect 441876 510992 445390 511048
rect 445446 510992 445451 511048
rect 441876 510990 445451 510992
rect 445385 510987 445451 510990
rect 444741 510506 444807 510509
rect 441876 510504 444807 510506
rect 441876 510448 444746 510504
rect 444802 510448 444807 510504
rect 441876 510446 444807 510448
rect 444741 510443 444807 510446
rect 370957 510098 371023 510101
rect 516133 510098 516199 510101
rect 369932 510096 371023 510098
rect 369932 510040 370962 510096
rect 371018 510040 371023 510096
rect 369932 510038 371023 510040
rect 513820 510096 516199 510098
rect 513820 510040 516138 510096
rect 516194 510040 516199 510096
rect 513820 510038 516199 510040
rect 370957 510035 371023 510038
rect 516133 510035 516199 510038
rect 445661 509962 445727 509965
rect 441876 509960 445727 509962
rect 441876 509904 445666 509960
rect 445722 509904 445727 509960
rect 441876 509902 445727 509904
rect 445661 509899 445727 509902
rect 369945 509418 370011 509421
rect 445569 509418 445635 509421
rect 369902 509416 370011 509418
rect 369902 509360 369950 509416
rect 370006 509360 370011 509416
rect 369902 509355 370011 509360
rect 441876 509416 445635 509418
rect 441876 509360 445574 509416
rect 445630 509360 445635 509416
rect 441876 509358 445635 509360
rect 445569 509355 445635 509358
rect 369902 508844 369962 509355
rect 445569 508874 445635 508877
rect 516133 508874 516199 508877
rect 441876 508872 445635 508874
rect 441876 508816 445574 508872
rect 445630 508816 445635 508872
rect 441876 508814 445635 508816
rect 513820 508872 516199 508874
rect 513820 508816 516138 508872
rect 516194 508816 516199 508872
rect 513820 508814 516199 508816
rect 445569 508811 445635 508814
rect 516133 508811 516199 508814
rect 445661 508330 445727 508333
rect 441876 508328 445727 508330
rect 441876 508272 445666 508328
rect 445722 508272 445727 508328
rect 441876 508270 445727 508272
rect 445661 508267 445727 508270
rect 516409 507786 516475 507789
rect 513820 507784 516475 507786
rect 369534 507517 369594 507756
rect 369485 507512 369594 507517
rect 369485 507456 369490 507512
rect 369546 507456 369594 507512
rect 369485 507454 369594 507456
rect 369485 507451 369551 507454
rect 441662 507381 441722 507756
rect 513820 507728 516414 507784
rect 516470 507728 516475 507784
rect 513820 507726 516475 507728
rect 516409 507723 516475 507726
rect 441662 507376 441771 507381
rect 441662 507320 441710 507376
rect 441766 507320 441771 507376
rect 441662 507318 441771 507320
rect 441705 507315 441771 507318
rect 445569 507242 445635 507245
rect 441876 507240 445635 507242
rect 441876 507184 445574 507240
rect 445630 507184 445635 507240
rect 441876 507182 445635 507184
rect 445569 507179 445635 507182
rect 445661 506698 445727 506701
rect 441876 506696 445727 506698
rect 441876 506640 445666 506696
rect 445722 506640 445727 506696
rect 441876 506638 445727 506640
rect 445661 506635 445727 506638
rect 370957 506562 371023 506565
rect 516133 506562 516199 506565
rect 369932 506560 371023 506562
rect 369932 506504 370962 506560
rect 371018 506504 371023 506560
rect 369932 506502 371023 506504
rect 513820 506560 516199 506562
rect 513820 506504 516138 506560
rect 516194 506504 516199 506560
rect 513820 506502 516199 506504
rect 370957 506499 371023 506502
rect 516133 506499 516199 506502
rect 445661 506154 445727 506157
rect 441876 506152 445727 506154
rect 441876 506096 445666 506152
rect 445722 506096 445727 506152
rect 441876 506094 445727 506096
rect 445661 506091 445727 506094
rect 445569 505610 445635 505613
rect 441876 505608 445635 505610
rect 441876 505552 445574 505608
rect 445630 505552 445635 505608
rect 441876 505550 445635 505552
rect 445569 505547 445635 505550
rect 516961 505474 517027 505477
rect 513820 505472 517027 505474
rect 369902 504930 369962 505444
rect 513820 505416 516966 505472
rect 517022 505416 517027 505472
rect 513820 505414 517027 505416
rect 516961 505411 517027 505414
rect 370037 504930 370103 504933
rect 369902 504928 370103 504930
rect 369902 504872 370042 504928
rect 370098 504872 370103 504928
rect 369902 504870 370103 504872
rect 370037 504867 370103 504870
rect 441662 504661 441722 505036
rect 441613 504656 441722 504661
rect 441613 504600 441618 504656
rect 441674 504600 441722 504656
rect 441613 504598 441722 504600
rect 441613 504595 441679 504598
rect 445661 504522 445727 504525
rect 441876 504520 445727 504522
rect 441876 504464 445666 504520
rect 445722 504464 445727 504520
rect 441876 504462 445727 504464
rect 445661 504459 445727 504462
rect 370957 504250 371023 504253
rect 516133 504250 516199 504253
rect 369932 504248 371023 504250
rect 369932 504192 370962 504248
rect 371018 504192 371023 504248
rect 369932 504190 371023 504192
rect 513820 504248 516199 504250
rect 513820 504192 516138 504248
rect 516194 504192 516199 504248
rect 513820 504190 516199 504192
rect 370957 504187 371023 504190
rect 516133 504187 516199 504190
rect 445293 504114 445359 504117
rect 441876 504112 445359 504114
rect 441876 504056 445298 504112
rect 445354 504056 445359 504112
rect 441876 504054 445359 504056
rect 445293 504051 445359 504054
rect 445109 503570 445175 503573
rect 441876 503568 445175 503570
rect 441876 503512 445114 503568
rect 445170 503512 445175 503568
rect 441876 503510 445175 503512
rect 445109 503507 445175 503510
rect 370957 503162 371023 503165
rect 516317 503162 516383 503165
rect 369932 503160 371023 503162
rect 369932 503104 370962 503160
rect 371018 503104 371023 503160
rect 369932 503102 371023 503104
rect 513820 503160 516383 503162
rect 513820 503104 516322 503160
rect 516378 503104 516383 503160
rect 513820 503102 516383 503104
rect 370957 503099 371023 503102
rect 516317 503099 516383 503102
rect 445017 503026 445083 503029
rect 441876 503024 445083 503026
rect 441876 502968 445022 503024
rect 445078 502968 445083 503024
rect 441876 502966 445083 502968
rect 445017 502963 445083 502966
rect 445201 502482 445267 502485
rect 441876 502480 445267 502482
rect 441876 502424 445206 502480
rect 445262 502424 445267 502480
rect 441876 502422 445267 502424
rect 445201 502419 445267 502422
rect 370129 501938 370195 501941
rect 445477 501938 445543 501941
rect 516869 501938 516935 501941
rect 369932 501936 370195 501938
rect -960 501802 480 501892
rect 369932 501880 370134 501936
rect 370190 501880 370195 501936
rect 369932 501878 370195 501880
rect 441876 501936 445543 501938
rect 441876 501880 445482 501936
rect 445538 501880 445543 501936
rect 441876 501878 445543 501880
rect 513820 501936 516935 501938
rect 513820 501880 516874 501936
rect 516930 501880 516935 501936
rect 513820 501878 516935 501880
rect 370129 501875 370195 501878
rect 445477 501875 445543 501878
rect 516869 501875 516935 501878
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 445293 501394 445359 501397
rect 441876 501392 445359 501394
rect 441876 501336 445298 501392
rect 445354 501336 445359 501392
rect 441876 501334 445359 501336
rect 445293 501331 445359 501334
rect 372521 500850 372587 500853
rect 444782 500850 444788 500852
rect 369932 500848 372587 500850
rect 369932 500792 372526 500848
rect 372582 500792 372587 500848
rect 369932 500790 372587 500792
rect 441876 500790 444788 500850
rect 372521 500787 372587 500790
rect 444782 500788 444788 500790
rect 444852 500788 444858 500852
rect 516133 500850 516199 500853
rect 513820 500848 516199 500850
rect 513820 500792 516138 500848
rect 516194 500792 516199 500848
rect 513820 500790 516199 500792
rect 516133 500787 516199 500790
rect 444414 500306 444420 500308
rect 441876 500246 444420 500306
rect 444414 500244 444420 500246
rect 444484 500306 444490 500308
rect 445569 500306 445635 500309
rect 444484 500304 445635 500306
rect 444484 500248 445574 500304
rect 445630 500248 445635 500304
rect 444484 500246 445635 500248
rect 444484 500244 444490 500246
rect 445569 500243 445635 500246
rect 445661 499762 445727 499765
rect 441876 499760 445727 499762
rect 441876 499704 445666 499760
rect 445722 499704 445727 499760
rect 441876 499702 445727 499704
rect 445661 499699 445727 499702
rect 370957 499626 371023 499629
rect 516133 499626 516199 499629
rect 369932 499624 371023 499626
rect 369932 499568 370962 499624
rect 371018 499568 371023 499624
rect 369932 499566 371023 499568
rect 513820 499624 516199 499626
rect 513820 499568 516138 499624
rect 516194 499568 516199 499624
rect 513820 499566 516199 499568
rect 370957 499563 371023 499566
rect 516133 499563 516199 499566
rect 445569 499218 445635 499221
rect 441876 499216 445635 499218
rect 441876 499160 445574 499216
rect 445630 499160 445635 499216
rect 441876 499158 445635 499160
rect 445569 499155 445635 499158
rect 444649 498674 444715 498677
rect 441876 498672 444715 498674
rect 441876 498616 444654 498672
rect 444710 498616 444715 498672
rect 441876 498614 444715 498616
rect 444649 498611 444715 498614
rect 370957 498538 371023 498541
rect 516133 498538 516199 498541
rect 369932 498536 371023 498538
rect 369932 498480 370962 498536
rect 371018 498480 371023 498536
rect 369932 498478 371023 498480
rect 513820 498536 516199 498538
rect 513820 498480 516138 498536
rect 516194 498480 516199 498536
rect 513820 498478 516199 498480
rect 370957 498475 371023 498478
rect 516133 498475 516199 498478
rect 445477 498130 445543 498133
rect 441876 498128 445543 498130
rect 441876 498072 445482 498128
rect 445538 498072 445543 498128
rect 441876 498070 445543 498072
rect 445477 498067 445543 498070
rect 583520 497844 584960 498084
rect 445753 497586 445819 497589
rect 441876 497584 445819 497586
rect 441876 497528 445758 497584
rect 445814 497528 445819 497584
rect 441876 497526 445819 497528
rect 445753 497523 445819 497526
rect 370221 497314 370287 497317
rect 516133 497314 516199 497317
rect 369932 497312 370287 497314
rect 369932 497256 370226 497312
rect 370282 497256 370287 497312
rect 369932 497254 370287 497256
rect 513820 497312 516199 497314
rect 513820 497256 516138 497312
rect 516194 497256 516199 497312
rect 513820 497254 516199 497256
rect 370221 497251 370287 497254
rect 516133 497251 516199 497254
rect 445569 497042 445635 497045
rect 441876 497040 445635 497042
rect 441876 496984 445574 497040
rect 445630 496984 445635 497040
rect 441876 496982 445635 496984
rect 445569 496979 445635 496982
rect 442993 496498 443059 496501
rect 443821 496498 443887 496501
rect 441876 496496 443887 496498
rect 441876 496440 442998 496496
rect 443054 496440 443826 496496
rect 443882 496440 443887 496496
rect 441876 496438 443887 496440
rect 442993 496435 443059 496438
rect 443821 496435 443887 496438
rect 370313 496226 370379 496229
rect 370681 496226 370747 496229
rect 516225 496226 516291 496229
rect 369932 496224 370747 496226
rect 369932 496168 370318 496224
rect 370374 496168 370686 496224
rect 370742 496168 370747 496224
rect 369932 496166 370747 496168
rect 513820 496224 516291 496226
rect 513820 496168 516230 496224
rect 516286 496168 516291 496224
rect 513820 496166 516291 496168
rect 370313 496163 370379 496166
rect 370681 496163 370747 496166
rect 516225 496163 516291 496166
rect 445845 495954 445911 495957
rect 441876 495952 445911 495954
rect 441876 495896 445850 495952
rect 445906 495896 445911 495952
rect 441876 495894 445911 495896
rect 445845 495891 445911 495894
rect 443085 495410 443151 495413
rect 443637 495410 443703 495413
rect 441876 495408 443703 495410
rect 441876 495352 443090 495408
rect 443146 495352 443642 495408
rect 443698 495352 443703 495408
rect 441876 495350 443703 495352
rect 443085 495347 443151 495350
rect 443637 495347 443703 495350
rect 370957 495002 371023 495005
rect 516869 495002 516935 495005
rect 517421 495002 517487 495005
rect 369932 495000 371023 495002
rect 369932 494944 370962 495000
rect 371018 494944 371023 495000
rect 369932 494942 371023 494944
rect 513820 495000 517487 495002
rect 513820 494944 516874 495000
rect 516930 494944 517426 495000
rect 517482 494944 517487 495000
rect 513820 494942 517487 494944
rect 370957 494939 371023 494942
rect 516869 494939 516935 494942
rect 517421 494939 517487 494942
rect 442901 494866 442967 494869
rect 441876 494864 442967 494866
rect 441876 494808 442906 494864
rect 442962 494808 442967 494864
rect 441876 494806 442967 494808
rect 442901 494803 442967 494806
rect 445293 494322 445359 494325
rect 441876 494320 445359 494322
rect 441876 494264 445298 494320
rect 445354 494264 445359 494320
rect 441876 494262 445359 494264
rect 445293 494259 445359 494262
rect 370957 493914 371023 493917
rect 442993 493914 443059 493917
rect 516317 493914 516383 493917
rect 517237 493914 517303 493917
rect 369932 493912 371023 493914
rect 369932 493856 370962 493912
rect 371018 493856 371023 493912
rect 369932 493854 371023 493856
rect 441876 493912 443059 493914
rect 441876 493856 442998 493912
rect 443054 493856 443059 493912
rect 441876 493854 443059 493856
rect 513820 493912 517303 493914
rect 513820 493856 516322 493912
rect 516378 493856 517242 493912
rect 517298 493856 517303 493912
rect 513820 493854 517303 493856
rect 370957 493851 371023 493854
rect 442993 493851 443059 493854
rect 516317 493851 516383 493854
rect 517237 493851 517303 493854
rect 445293 493370 445359 493373
rect 441876 493368 445359 493370
rect 441876 493312 445298 493368
rect 445354 493312 445359 493368
rect 441876 493310 445359 493312
rect 445293 493307 445359 493310
rect 444649 492826 444715 492829
rect 441876 492824 444715 492826
rect 441876 492768 444654 492824
rect 444710 492768 444715 492824
rect 441876 492766 444715 492768
rect 444649 492763 444715 492766
rect 370773 492690 370839 492693
rect 516225 492690 516291 492693
rect 369932 492688 370839 492690
rect 369932 492632 370778 492688
rect 370834 492632 370839 492688
rect 369932 492630 370839 492632
rect 513820 492688 516291 492690
rect 513820 492632 516230 492688
rect 516286 492632 516291 492688
rect 513820 492630 516291 492632
rect 370773 492627 370839 492630
rect 516225 492627 516291 492630
rect 441797 492554 441863 492557
rect 441797 492552 441906 492554
rect 441797 492496 441802 492552
rect 441858 492496 441906 492552
rect 441797 492491 441906 492496
rect 441846 492282 441906 492491
rect 442533 492282 442599 492285
rect 441846 492280 442599 492282
rect 441846 492252 442538 492280
rect 441876 492224 442538 492252
rect 442594 492224 442599 492280
rect 441876 492222 442599 492224
rect 442533 492219 442599 492222
rect 443545 491738 443611 491741
rect 441876 491736 443611 491738
rect 441876 491680 443550 491736
rect 443606 491680 443611 491736
rect 441876 491678 443611 491680
rect 443545 491675 443611 491678
rect 370865 491602 370931 491605
rect 516133 491602 516199 491605
rect 369932 491600 370931 491602
rect 369932 491544 370870 491600
rect 370926 491544 370931 491600
rect 369932 491542 370931 491544
rect 513820 491600 516199 491602
rect 513820 491544 516138 491600
rect 516194 491544 516199 491600
rect 513820 491542 516199 491544
rect 370865 491539 370931 491542
rect 516133 491539 516199 491542
rect 445293 491194 445359 491197
rect 441876 491192 445359 491194
rect 441876 491136 445298 491192
rect 445354 491136 445359 491192
rect 441876 491134 445359 491136
rect 445293 491131 445359 491134
rect 443177 490650 443243 490653
rect 441876 490648 443243 490650
rect 441876 490592 443182 490648
rect 443238 490592 443243 490648
rect 441876 490590 443243 490592
rect 443177 490587 443243 490590
rect 370957 490378 371023 490381
rect 516133 490378 516199 490381
rect 369932 490376 371023 490378
rect 369932 490320 370962 490376
rect 371018 490320 371023 490376
rect 369932 490318 371023 490320
rect 513820 490376 516199 490378
rect 513820 490320 516138 490376
rect 516194 490320 516199 490376
rect 513820 490318 516199 490320
rect 370957 490315 371023 490318
rect 516133 490315 516199 490318
rect 443913 490106 443979 490109
rect 441876 490104 443979 490106
rect 441876 490048 443918 490104
rect 443974 490048 443979 490104
rect 441876 490046 443979 490048
rect 443913 490043 443979 490046
rect 441889 489698 441955 489701
rect 441846 489696 441955 489698
rect 441846 489640 441894 489696
rect 441950 489640 441955 489696
rect 441846 489635 441955 489640
rect 441846 489532 441906 489635
rect 370405 489290 370471 489293
rect 516685 489290 516751 489293
rect 369932 489288 370471 489290
rect 369932 489232 370410 489288
rect 370466 489232 370471 489288
rect 513452 489288 516751 489290
rect 513452 489260 516690 489288
rect 369932 489230 370471 489232
rect 370405 489227 370471 489230
rect 513422 489232 516690 489260
rect 516746 489232 516751 489288
rect 513422 489230 516751 489232
rect 443453 489018 443519 489021
rect 441876 489016 443519 489018
rect 441876 488960 443458 489016
rect 443514 488960 443519 489016
rect 441876 488958 443519 488960
rect 443453 488955 443519 488958
rect -960 488596 480 488836
rect 513422 488749 513482 489230
rect 516685 489227 516751 489230
rect 513422 488744 513531 488749
rect 513422 488688 513470 488744
rect 513526 488688 513531 488744
rect 513422 488686 513531 488688
rect 513465 488683 513531 488686
rect 445477 488474 445543 488477
rect 441876 488472 445543 488474
rect 441876 488416 445482 488472
rect 445538 488416 445543 488472
rect 441876 488414 445543 488416
rect 445477 488411 445543 488414
rect 369761 488202 369827 488205
rect 369718 488200 369827 488202
rect 369718 488144 369766 488200
rect 369822 488144 369827 488200
rect 369718 488139 369827 488144
rect 369718 488036 369778 488139
rect 517237 488066 517303 488069
rect 513452 488064 517303 488066
rect 513452 488036 517242 488064
rect 513422 488008 517242 488036
rect 517298 488008 517303 488064
rect 513422 488006 517303 488008
rect 444649 487930 444715 487933
rect 441876 487928 444715 487930
rect 441876 487872 444654 487928
rect 444710 487872 444715 487928
rect 441876 487870 444715 487872
rect 444649 487867 444715 487870
rect 513422 487525 513482 488006
rect 517237 488003 517303 488006
rect 513373 487520 513482 487525
rect 513373 487464 513378 487520
rect 513434 487464 513482 487520
rect 513373 487462 513482 487464
rect 513373 487459 513439 487462
rect 445293 487386 445359 487389
rect 441876 487384 445359 487386
rect 441876 487328 445298 487384
rect 445354 487328 445359 487384
rect 441876 487326 445359 487328
rect 445293 487323 445359 487326
rect 372521 486978 372587 486981
rect 441981 486978 442047 486981
rect 516133 486978 516199 486981
rect 369932 486976 372587 486978
rect 369932 486920 372526 486976
rect 372582 486920 372587 486976
rect 369932 486918 372587 486920
rect 372521 486915 372587 486918
rect 441846 486976 442047 486978
rect 441846 486920 441986 486976
rect 442042 486920 442047 486976
rect 441846 486918 442047 486920
rect 513820 486976 516199 486978
rect 513820 486920 516138 486976
rect 516194 486920 516199 486976
rect 513820 486918 516199 486920
rect 441846 486434 441906 486918
rect 441981 486915 442047 486918
rect 516133 486915 516199 486918
rect 443269 486434 443335 486437
rect 441846 486432 443335 486434
rect 441846 486376 443274 486432
rect 443330 486376 443335 486432
rect 441846 486374 443335 486376
rect 443269 486371 443335 486374
rect 445477 486298 445543 486301
rect 441876 486296 445543 486298
rect 441876 486240 445482 486296
rect 445538 486240 445543 486296
rect 441876 486238 445543 486240
rect 445477 486235 445543 486238
rect 370957 485754 371023 485757
rect 442625 485754 442691 485757
rect 445109 485754 445175 485757
rect 516133 485754 516199 485757
rect 369932 485752 371023 485754
rect 369932 485696 370962 485752
rect 371018 485696 371023 485752
rect 369932 485694 371023 485696
rect 441876 485752 445175 485754
rect 441876 485696 442630 485752
rect 442686 485696 445114 485752
rect 445170 485696 445175 485752
rect 513820 485752 516199 485754
rect 513820 485724 516138 485752
rect 441876 485694 445175 485696
rect 370957 485691 371023 485694
rect 442625 485691 442691 485694
rect 445109 485691 445175 485694
rect 513790 485696 516138 485724
rect 516194 485696 516199 485752
rect 513790 485694 516199 485696
rect 513790 485213 513850 485694
rect 516133 485691 516199 485694
rect 442073 485210 442139 485213
rect 441876 485208 442139 485210
rect 441876 485180 442078 485208
rect 441846 485152 442078 485180
rect 442134 485152 442139 485208
rect 441846 485150 442139 485152
rect 441846 484802 441906 485150
rect 442073 485147 442139 485150
rect 513741 485208 513850 485213
rect 513741 485152 513746 485208
rect 513802 485152 513850 485208
rect 513741 485150 513850 485152
rect 513741 485147 513807 485150
rect 443361 484802 443427 484805
rect 441846 484800 443427 484802
rect 441846 484744 443366 484800
rect 443422 484744 443427 484800
rect 441846 484742 443427 484744
rect 443361 484739 443427 484742
rect 370497 484666 370563 484669
rect 445477 484666 445543 484669
rect 517605 484666 517671 484669
rect 369932 484664 370563 484666
rect 369932 484608 370502 484664
rect 370558 484608 370563 484664
rect 369932 484606 370563 484608
rect 441876 484664 445543 484666
rect 441876 484608 445482 484664
rect 445538 484608 445543 484664
rect 441876 484606 445543 484608
rect 513820 484664 517671 484666
rect 513820 484608 517610 484664
rect 517666 484608 517671 484664
rect 513820 484606 517671 484608
rect 370497 484603 370563 484606
rect 445477 484603 445543 484606
rect 517605 484603 517671 484606
rect 582465 484666 582531 484669
rect 583520 484666 584960 484756
rect 582465 484664 584960 484666
rect 582465 484608 582470 484664
rect 582526 484608 584960 484664
rect 582465 484606 584960 484608
rect 582465 484603 582531 484606
rect 583520 484516 584960 484606
rect 444649 484258 444715 484261
rect 441876 484256 444715 484258
rect 441876 484200 444654 484256
rect 444710 484200 444715 484256
rect 441876 484198 444715 484200
rect 444649 484195 444715 484198
rect 365161 484122 365227 484125
rect 365294 484122 365300 484124
rect 365161 484120 365300 484122
rect 365161 484064 365166 484120
rect 365222 484064 365300 484120
rect 365161 484062 365300 484064
rect 365161 484059 365227 484062
rect 365294 484060 365300 484062
rect 365364 484060 365370 484124
rect 435173 483988 435239 483989
rect 436737 483988 436803 483989
rect 435173 483984 435220 483988
rect 435284 483986 435290 483988
rect 436686 483986 436692 483988
rect 435173 483928 435178 483984
rect 435173 483924 435220 483928
rect 435284 483926 435330 483986
rect 436646 483926 436692 483986
rect 436756 483984 436803 483988
rect 436798 483928 436803 483984
rect 435284 483924 435290 483926
rect 436686 483924 436692 483926
rect 436756 483924 436803 483928
rect 435173 483923 435239 483924
rect 436737 483923 436803 483924
rect 365294 482836 365300 482900
rect 365364 482898 365370 482900
rect 371141 482898 371207 482901
rect 365364 482896 371207 482898
rect 365364 482840 371146 482896
rect 371202 482840 371207 482896
rect 365364 482838 371207 482840
rect 365364 482836 365370 482838
rect 371141 482835 371207 482838
rect 361614 482156 361620 482220
rect 361684 482218 361690 482220
rect 362718 482218 362724 482220
rect 361684 482158 362724 482218
rect 361684 482156 361690 482158
rect 362718 482156 362724 482158
rect 362788 482218 362794 482220
rect 362861 482218 362927 482221
rect 362788 482216 362927 482218
rect 362788 482160 362866 482216
rect 362922 482160 362927 482216
rect 362788 482158 362927 482160
rect 362788 482156 362794 482158
rect 362861 482155 362927 482158
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect 371325 441826 371391 441829
rect 369902 441824 371391 441826
rect 369902 441768 371330 441824
rect 371386 441768 371391 441824
rect 369902 441766 371391 441768
rect 369902 441660 369962 441766
rect 371325 441763 371391 441766
rect 517053 441690 517119 441693
rect 513820 441688 517119 441690
rect 513820 441632 517058 441688
rect 517114 441632 517119 441688
rect 513820 441630 517119 441632
rect 517053 441627 517119 441630
rect 445109 441418 445175 441421
rect 441876 441416 445175 441418
rect 441876 441360 445114 441416
rect 445170 441360 445175 441416
rect 441876 441358 445175 441360
rect 445109 441355 445175 441358
rect 371233 441146 371299 441149
rect 517329 441146 517395 441149
rect 369932 441144 371299 441146
rect 369932 441088 371238 441144
rect 371294 441088 371299 441144
rect 369932 441086 371299 441088
rect 513820 441144 517395 441146
rect 513820 441088 517334 441144
rect 517390 441088 517395 441144
rect 513820 441086 517395 441088
rect 371233 441083 371299 441086
rect 517329 441083 517395 441086
rect 371417 440602 371483 440605
rect 516133 440602 516199 440605
rect 369932 440600 371483 440602
rect 369932 440544 371422 440600
rect 371478 440544 371483 440600
rect 513820 440600 516199 440602
rect 513820 440572 516138 440600
rect 369932 440542 371483 440544
rect 371417 440539 371483 440542
rect 513790 440544 516138 440572
rect 516194 440544 516199 440600
rect 513790 440542 516199 440544
rect 371233 440466 371299 440469
rect 371877 440466 371943 440469
rect 371233 440464 371943 440466
rect 371233 440408 371238 440464
rect 371294 440408 371882 440464
rect 371938 440408 371943 440464
rect 371233 440406 371943 440408
rect 371233 440403 371299 440406
rect 371877 440403 371943 440406
rect 513790 440333 513850 440542
rect 516133 440539 516199 440542
rect 445569 440330 445635 440333
rect 441876 440328 445635 440330
rect 441876 440272 445574 440328
rect 445630 440272 445635 440328
rect 441876 440270 445635 440272
rect 445569 440267 445635 440270
rect 513741 440328 513850 440333
rect 513741 440272 513746 440328
rect 513802 440272 513850 440328
rect 513741 440270 513850 440272
rect 513741 440267 513807 440270
rect 371182 440058 371188 440060
rect 369932 439998 371188 440058
rect 371182 439996 371188 439998
rect 371252 439996 371258 440060
rect 517237 440058 517303 440061
rect 513820 440056 517303 440058
rect 513820 440000 517242 440056
rect 517298 440000 517303 440056
rect 513820 439998 517303 440000
rect 517237 439995 517303 439998
rect 371366 439514 371372 439516
rect 369932 439454 371372 439514
rect 371366 439452 371372 439454
rect 371436 439452 371442 439516
rect 516174 439514 516180 439516
rect 513820 439454 516180 439514
rect 516174 439452 516180 439454
rect 516244 439452 516250 439516
rect 371182 439044 371188 439108
rect 371252 439106 371258 439108
rect 372470 439106 372476 439108
rect 371252 439046 372476 439106
rect 371252 439044 371258 439046
rect 372470 439044 372476 439046
rect 372540 439044 372546 439108
rect 443821 439106 443887 439109
rect 444189 439106 444255 439109
rect 441876 439104 444255 439106
rect 441876 439048 443826 439104
rect 443882 439048 444194 439104
rect 444250 439048 444255 439104
rect 441876 439046 444255 439048
rect 443821 439043 443887 439046
rect 444189 439043 444255 439046
rect 371182 438970 371188 438972
rect 369932 438910 371188 438970
rect 371182 438908 371188 438910
rect 371252 438970 371258 438972
rect 371550 438970 371556 438972
rect 371252 438910 371556 438970
rect 371252 438908 371258 438910
rect 371550 438908 371556 438910
rect 371620 438908 371626 438972
rect 516133 438970 516199 438973
rect 513820 438968 516199 438970
rect 513820 438912 516138 438968
rect 516194 438912 516199 438968
rect 513820 438910 516199 438912
rect 516133 438907 516199 438910
rect 371785 438426 371851 438429
rect 516225 438426 516291 438429
rect 369932 438424 371851 438426
rect 369932 438368 371790 438424
rect 371846 438368 371851 438424
rect 369932 438366 371851 438368
rect 513820 438424 516291 438426
rect 513820 438368 516230 438424
rect 516286 438368 516291 438424
rect 513820 438366 516291 438368
rect 371785 438363 371851 438366
rect 516225 438363 516291 438366
rect 444649 438018 444715 438021
rect 441876 438016 444715 438018
rect 441876 437960 444654 438016
rect 444710 437960 444715 438016
rect 441876 437958 444715 437960
rect 444649 437955 444715 437958
rect 371601 437882 371667 437885
rect 516133 437882 516199 437885
rect 369932 437880 371667 437882
rect 369932 437824 371606 437880
rect 371662 437824 371667 437880
rect 369932 437822 371667 437824
rect 513820 437880 516199 437882
rect 513820 437824 516138 437880
rect 516194 437824 516199 437880
rect 513820 437822 516199 437824
rect 371601 437819 371667 437822
rect 516133 437819 516199 437822
rect 371693 437338 371759 437341
rect 516225 437338 516291 437341
rect 369932 437336 371759 437338
rect 369932 437280 371698 437336
rect 371754 437280 371759 437336
rect 369932 437278 371759 437280
rect 513820 437336 516291 437338
rect 513820 437280 516230 437336
rect 516286 437280 516291 437336
rect 513820 437278 516291 437280
rect 371693 437275 371759 437278
rect 516225 437275 516291 437278
rect 371601 436794 371667 436797
rect 444373 436794 444439 436797
rect 516501 436794 516567 436797
rect 369932 436792 371667 436794
rect -960 436508 480 436748
rect 369932 436736 371606 436792
rect 371662 436736 371667 436792
rect 369932 436734 371667 436736
rect 441876 436792 444439 436794
rect 441876 436736 444378 436792
rect 444434 436736 444439 436792
rect 441876 436734 444439 436736
rect 513820 436792 516567 436794
rect 513820 436736 516506 436792
rect 516562 436736 516567 436792
rect 513820 436734 516567 436736
rect 371601 436731 371667 436734
rect 444373 436731 444439 436734
rect 516501 436731 516567 436734
rect 371785 436250 371851 436253
rect 516133 436250 516199 436253
rect 369932 436248 371851 436250
rect 369932 436192 371790 436248
rect 371846 436192 371851 436248
rect 369932 436190 371851 436192
rect 513820 436248 516199 436250
rect 513820 436192 516138 436248
rect 516194 436192 516199 436248
rect 513820 436190 516199 436192
rect 371785 436187 371851 436190
rect 516133 436187 516199 436190
rect 371601 435706 371667 435709
rect 442441 435706 442507 435709
rect 516225 435706 516291 435709
rect 369932 435704 371667 435706
rect 369932 435648 371606 435704
rect 371662 435648 371667 435704
rect 441876 435704 442507 435706
rect 441876 435676 442446 435704
rect 369932 435646 371667 435648
rect 371601 435643 371667 435646
rect 441846 435648 442446 435676
rect 442502 435648 442507 435704
rect 441846 435646 442507 435648
rect 513820 435704 516291 435706
rect 513820 435648 516230 435704
rect 516286 435648 516291 435704
rect 513820 435646 516291 435648
rect 441846 435573 441906 435646
rect 442441 435643 442507 435646
rect 516225 435643 516291 435646
rect 441797 435568 441906 435573
rect 441797 435512 441802 435568
rect 441858 435512 441906 435568
rect 441797 435510 441906 435512
rect 441797 435507 441863 435510
rect 371693 435162 371759 435165
rect 516133 435162 516199 435165
rect 369932 435160 371759 435162
rect 369932 435104 371698 435160
rect 371754 435104 371759 435160
rect 369932 435102 371759 435104
rect 513820 435160 516199 435162
rect 513820 435104 516138 435160
rect 516194 435104 516199 435160
rect 513820 435102 516199 435104
rect 371693 435099 371759 435102
rect 516133 435099 516199 435102
rect 371601 434618 371667 434621
rect 516501 434618 516567 434621
rect 369932 434616 371667 434618
rect 369932 434560 371606 434616
rect 371662 434560 371667 434616
rect 369932 434558 371667 434560
rect 513820 434616 516567 434618
rect 513820 434560 516506 434616
rect 516562 434560 516567 434616
rect 513820 434558 516567 434560
rect 371601 434555 371667 434558
rect 516501 434555 516567 434558
rect 444465 434482 444531 434485
rect 441876 434480 444531 434482
rect 441876 434424 444470 434480
rect 444526 434424 444531 434480
rect 441876 434422 444531 434424
rect 444465 434419 444531 434422
rect 371693 434074 371759 434077
rect 516225 434074 516291 434077
rect 369932 434072 371759 434074
rect 369932 434016 371698 434072
rect 371754 434016 371759 434072
rect 369932 434014 371759 434016
rect 513820 434072 516291 434074
rect 513820 434016 516230 434072
rect 516286 434016 516291 434072
rect 513820 434014 516291 434016
rect 371693 434011 371759 434014
rect 516225 434011 516291 434014
rect 371785 433530 371851 433533
rect 516133 433530 516199 433533
rect 369932 433528 371851 433530
rect 369932 433472 371790 433528
rect 371846 433472 371851 433528
rect 369932 433470 371851 433472
rect 513820 433528 516199 433530
rect 513820 433472 516138 433528
rect 516194 433472 516199 433528
rect 513820 433470 516199 433472
rect 371785 433467 371851 433470
rect 516133 433467 516199 433470
rect 442993 433394 443059 433397
rect 441876 433392 443059 433394
rect 441876 433336 442998 433392
rect 443054 433336 443059 433392
rect 441876 433334 443059 433336
rect 442993 433331 443059 433334
rect 371693 432986 371759 432989
rect 516501 432986 516567 432989
rect 369932 432984 371759 432986
rect 369932 432928 371698 432984
rect 371754 432928 371759 432984
rect 369932 432926 371759 432928
rect 513820 432984 516567 432986
rect 513820 432928 516506 432984
rect 516562 432928 516567 432984
rect 513820 432926 516567 432928
rect 371693 432923 371759 432926
rect 516501 432923 516567 432926
rect 371601 432442 371667 432445
rect 516777 432442 516843 432445
rect 369932 432440 371667 432442
rect 369932 432384 371606 432440
rect 371662 432384 371667 432440
rect 369932 432382 371667 432384
rect 513820 432440 516843 432442
rect 513820 432384 516782 432440
rect 516838 432384 516843 432440
rect 513820 432382 516843 432384
rect 371601 432379 371667 432382
rect 516777 432379 516843 432382
rect 513465 432306 513531 432309
rect 513422 432304 513531 432306
rect 513422 432248 513470 432304
rect 513526 432248 513531 432304
rect 513422 432243 513531 432248
rect 444465 432170 444531 432173
rect 441876 432168 444531 432170
rect 441876 432112 444470 432168
rect 444526 432112 444531 432168
rect 441876 432110 444531 432112
rect 444465 432107 444531 432110
rect 371601 432034 371667 432037
rect 369932 432032 371667 432034
rect 369932 431976 371606 432032
rect 371662 431976 371667 432032
rect 513422 432004 513482 432243
rect 516225 432034 516291 432037
rect 516869 432034 516935 432037
rect 516225 432032 516935 432034
rect 369932 431974 371667 431976
rect 371601 431971 371667 431974
rect 516225 431976 516230 432032
rect 516286 431976 516874 432032
rect 516930 431976 516935 432032
rect 516225 431974 516935 431976
rect 516225 431971 516291 431974
rect 516869 431971 516935 431974
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 371693 431490 371759 431493
rect 516225 431490 516291 431493
rect 369932 431488 371759 431490
rect 369932 431432 371698 431488
rect 371754 431432 371759 431488
rect 369932 431430 371759 431432
rect 513820 431488 516291 431490
rect 513820 431432 516230 431488
rect 516286 431432 516291 431488
rect 583520 431476 584960 431566
rect 513820 431430 516291 431432
rect 371693 431427 371759 431430
rect 516225 431427 516291 431430
rect 443085 431082 443151 431085
rect 441876 431080 443151 431082
rect 441876 431024 443090 431080
rect 443146 431024 443151 431080
rect 441876 431022 443151 431024
rect 443085 431019 443151 431022
rect 371509 430946 371575 430949
rect 516409 430946 516475 430949
rect 369932 430944 371575 430946
rect 369932 430888 371514 430944
rect 371570 430888 371575 430944
rect 369932 430886 371575 430888
rect 513820 430944 516475 430946
rect 513820 430888 516414 430944
rect 516470 430888 516475 430944
rect 513820 430886 516475 430888
rect 371509 430883 371575 430886
rect 516409 430883 516475 430886
rect 371693 430674 371759 430677
rect 371877 430674 371943 430677
rect 371693 430672 371943 430674
rect 371693 430616 371698 430672
rect 371754 430616 371882 430672
rect 371938 430616 371943 430672
rect 371693 430614 371943 430616
rect 371693 430611 371759 430614
rect 371877 430611 371943 430614
rect 513373 430674 513439 430677
rect 513373 430672 513482 430674
rect 513373 430616 513378 430672
rect 513434 430616 513482 430672
rect 513373 430611 513482 430616
rect 372153 430402 372219 430405
rect 369932 430400 372219 430402
rect 369932 430344 372158 430400
rect 372214 430344 372219 430400
rect 513422 430372 513482 430611
rect 369932 430342 372219 430344
rect 372153 430339 372219 430342
rect 371969 429858 372035 429861
rect 442533 429858 442599 429861
rect 516409 429858 516475 429861
rect 369932 429856 372035 429858
rect 369932 429800 371974 429856
rect 372030 429800 372035 429856
rect 441876 429856 442599 429858
rect 441876 429828 442538 429856
rect 369932 429798 372035 429800
rect 371969 429795 372035 429798
rect 441846 429800 442538 429828
rect 442594 429800 442599 429856
rect 441846 429798 442599 429800
rect 513820 429856 516475 429858
rect 513820 429800 516414 429856
rect 516470 429800 516475 429856
rect 513820 429798 516475 429800
rect 441846 429317 441906 429798
rect 442533 429795 442599 429798
rect 516409 429795 516475 429798
rect 372061 429314 372127 429317
rect 369932 429312 372127 429314
rect 369932 429256 372066 429312
rect 372122 429256 372127 429312
rect 369932 429254 372127 429256
rect 441846 429312 441955 429317
rect 516501 429314 516567 429317
rect 441846 429256 441894 429312
rect 441950 429256 441955 429312
rect 441846 429254 441955 429256
rect 513820 429312 516567 429314
rect 513820 429256 516506 429312
rect 516562 429256 516567 429312
rect 513820 429254 516567 429256
rect 372061 429251 372127 429254
rect 441889 429251 441955 429254
rect 516501 429251 516567 429254
rect 371918 428770 371924 428772
rect 369932 428710 371924 428770
rect 371918 428708 371924 428710
rect 371988 428770 371994 428772
rect 372245 428770 372311 428773
rect 442073 428770 442139 428773
rect 516409 428770 516475 428773
rect 371988 428768 372311 428770
rect 371988 428712 372250 428768
rect 372306 428712 372311 428768
rect 371988 428710 372311 428712
rect 441876 428768 442139 428770
rect 441876 428712 442078 428768
rect 442134 428712 442139 428768
rect 441876 428710 442139 428712
rect 513820 428768 516475 428770
rect 513820 428712 516414 428768
rect 516470 428712 516475 428768
rect 513820 428710 516475 428712
rect 371988 428708 371994 428710
rect 372245 428707 372311 428710
rect 442073 428707 442139 428710
rect 516409 428707 516475 428710
rect 371734 428226 371740 428228
rect 369932 428166 371740 428226
rect 371734 428164 371740 428166
rect 371804 428164 371810 428228
rect 516777 428226 516843 428229
rect 513820 428224 516843 428226
rect 513820 428168 516782 428224
rect 516838 428168 516843 428224
rect 513820 428166 516843 428168
rect 516777 428163 516843 428166
rect 516961 427682 517027 427685
rect 513820 427680 517027 427682
rect 369350 427412 369410 427652
rect 513820 427624 516966 427680
rect 517022 427624 517027 427680
rect 513820 427622 517027 427624
rect 516961 427619 517027 427622
rect 445937 427546 446003 427549
rect 441876 427544 446003 427546
rect 441876 427488 445942 427544
rect 445998 427488 446003 427544
rect 441876 427486 446003 427488
rect 445937 427483 446003 427486
rect 369342 427348 369348 427412
rect 369412 427410 369418 427412
rect 371233 427410 371299 427413
rect 369412 427408 371299 427410
rect 369412 427352 371238 427408
rect 371294 427352 371299 427408
rect 369412 427350 371299 427352
rect 369412 427348 369418 427350
rect 371233 427347 371299 427350
rect 371601 427138 371667 427141
rect 516685 427138 516751 427141
rect 369932 427136 371667 427138
rect 369932 427080 371606 427136
rect 371662 427080 371667 427136
rect 369932 427078 371667 427080
rect 513820 427136 516751 427138
rect 513820 427080 516690 427136
rect 516746 427080 516751 427136
rect 513820 427078 516751 427080
rect 371601 427075 371667 427078
rect 516685 427075 516751 427078
rect 371601 426594 371667 426597
rect 516133 426594 516199 426597
rect 369932 426592 371667 426594
rect 369932 426536 371606 426592
rect 371662 426536 371667 426592
rect 369932 426534 371667 426536
rect 513820 426592 516199 426594
rect 513820 426536 516138 426592
rect 516194 426536 516199 426592
rect 513820 426534 516199 426536
rect 371601 426531 371667 426534
rect 516133 426531 516199 426534
rect 445569 426458 445635 426461
rect 441876 426456 445635 426458
rect 441876 426400 445574 426456
rect 445630 426400 445635 426456
rect 441876 426398 445635 426400
rect 445569 426395 445635 426398
rect 371601 426050 371667 426053
rect 516317 426050 516383 426053
rect 369932 426048 371667 426050
rect 369932 425992 371606 426048
rect 371662 425992 371667 426048
rect 369932 425990 371667 425992
rect 513820 426048 516383 426050
rect 513820 425992 516322 426048
rect 516378 425992 516383 426048
rect 513820 425990 516383 425992
rect 371601 425987 371667 425990
rect 516317 425987 516383 425990
rect 369853 425914 369919 425917
rect 369853 425912 369962 425914
rect 369853 425856 369858 425912
rect 369914 425856 369962 425912
rect 369853 425851 369962 425856
rect 369902 425506 369962 425851
rect 371049 425506 371115 425509
rect 516777 425506 516843 425509
rect 369902 425504 371115 425506
rect 369902 425476 371054 425504
rect 369932 425448 371054 425476
rect 371110 425448 371115 425504
rect 369932 425446 371115 425448
rect 513820 425504 516843 425506
rect 513820 425448 516782 425504
rect 516838 425448 516843 425504
rect 513820 425446 516843 425448
rect 371049 425443 371115 425446
rect 516777 425443 516843 425446
rect 369485 425234 369551 425237
rect 443545 425234 443611 425237
rect 443913 425234 443979 425237
rect 369485 425232 369594 425234
rect 369485 425176 369490 425232
rect 369546 425176 369594 425232
rect 369485 425171 369594 425176
rect 441876 425232 443979 425234
rect 441876 425176 443550 425232
rect 443606 425176 443918 425232
rect 443974 425176 443979 425232
rect 441876 425174 443979 425176
rect 443545 425171 443611 425174
rect 443913 425171 443979 425174
rect 369534 424962 369594 425171
rect 371233 424962 371299 424965
rect 516133 424962 516199 424965
rect 369534 424960 371299 424962
rect 369534 424932 371238 424960
rect 369564 424904 371238 424932
rect 371294 424904 371299 424960
rect 369564 424902 371299 424904
rect 513820 424960 516199 424962
rect 513820 424904 516138 424960
rect 516194 424904 516199 424960
rect 513820 424902 516199 424904
rect 371233 424899 371299 424902
rect 516133 424899 516199 424902
rect 372613 424418 372679 424421
rect 516133 424418 516199 424421
rect 369932 424416 372679 424418
rect 369932 424360 372618 424416
rect 372674 424360 372679 424416
rect 369932 424358 372679 424360
rect 513820 424416 516199 424418
rect 513820 424360 516138 424416
rect 516194 424360 516199 424416
rect 513820 424358 516199 424360
rect 372613 424355 372679 424358
rect 516133 424355 516199 424358
rect 442349 424146 442415 424149
rect 441876 424144 442415 424146
rect 441876 424116 442354 424144
rect 441846 424088 442354 424116
rect 442410 424088 442415 424144
rect 441846 424086 442415 424088
rect 441846 424010 441906 424086
rect 442349 424083 442415 424086
rect 441981 424010 442047 424013
rect 441846 424008 442047 424010
rect 441846 423952 441986 424008
rect 442042 423952 442047 424008
rect 441846 423950 442047 423952
rect 441981 423947 442047 423950
rect 371601 423874 371667 423877
rect 516225 423874 516291 423877
rect 369932 423872 371667 423874
rect 369932 423816 371606 423872
rect 371662 423816 371667 423872
rect 369932 423814 371667 423816
rect 513820 423872 516291 423874
rect 513820 423816 516230 423872
rect 516286 423816 516291 423872
rect 513820 423814 516291 423816
rect 371601 423811 371667 423814
rect 516225 423811 516291 423814
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect 369945 423602 370011 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 369902 423600 370011 423602
rect 369902 423544 369950 423600
rect 370006 423544 370011 423600
rect 369902 423539 370011 423544
rect 369902 423330 369962 423539
rect 371141 423330 371207 423333
rect 516133 423330 516199 423333
rect 369902 423328 371207 423330
rect 369902 423300 371146 423328
rect 369932 423272 371146 423300
rect 371202 423272 371207 423328
rect 369932 423270 371207 423272
rect 513820 423328 516199 423330
rect 513820 423272 516138 423328
rect 516194 423272 516199 423328
rect 513820 423270 516199 423272
rect 371141 423267 371207 423270
rect 516133 423267 516199 423270
rect 369301 423194 369367 423197
rect 369301 423192 369410 423194
rect 369301 423136 369306 423192
rect 369362 423136 369410 423192
rect 369301 423131 369410 423136
rect 369350 422786 369410 423131
rect 442257 422922 442323 422925
rect 441876 422920 442323 422922
rect 441876 422864 442262 422920
rect 442318 422864 442323 422920
rect 441876 422862 442323 422864
rect 442257 422859 442323 422862
rect 516317 422786 516383 422789
rect 369350 422756 369932 422786
rect 513820 422784 516383 422786
rect 369380 422726 369962 422756
rect 513820 422728 516322 422784
rect 516378 422728 516383 422784
rect 513820 422726 516383 422728
rect 369902 422514 369962 422726
rect 516317 422723 516383 422726
rect 370405 422514 370471 422517
rect 369902 422512 370471 422514
rect 369902 422456 370410 422512
rect 370466 422456 370471 422512
rect 369902 422454 370471 422456
rect 370405 422451 370471 422454
rect 371969 422242 372035 422245
rect 516317 422242 516383 422245
rect 369932 422240 372035 422242
rect 369932 422184 371974 422240
rect 372030 422184 372035 422240
rect 369932 422182 372035 422184
rect 513820 422240 516383 422242
rect 513820 422184 516322 422240
rect 516378 422184 516383 422240
rect 513820 422182 516383 422184
rect 371969 422179 372035 422182
rect 516317 422179 516383 422182
rect 443821 421834 443887 421837
rect 516317 421834 516383 421837
rect 441876 421832 443887 421834
rect 369902 421698 369962 421804
rect 441876 421776 443826 421832
rect 443882 421776 443887 421832
rect 441876 421774 443887 421776
rect 513820 421832 516383 421834
rect 513820 421776 516322 421832
rect 516378 421776 516383 421832
rect 513820 421774 516383 421776
rect 443821 421771 443887 421774
rect 516317 421771 516383 421774
rect 370037 421698 370103 421701
rect 369902 421696 370103 421698
rect 369902 421640 370042 421696
rect 370098 421640 370103 421696
rect 369902 421638 370103 421640
rect 370037 421635 370103 421638
rect 373073 421290 373139 421293
rect 516317 421290 516383 421293
rect 369380 421288 373139 421290
rect 369380 421260 373078 421288
rect 369350 421232 373078 421260
rect 373134 421232 373139 421288
rect 369350 421230 373139 421232
rect 513820 421288 516383 421290
rect 513820 421232 516322 421288
rect 516378 421232 516383 421288
rect 513820 421230 516383 421232
rect 369350 421021 369410 421230
rect 373073 421227 373139 421230
rect 516317 421227 516383 421230
rect 369301 421016 369410 421021
rect 369301 420960 369306 421016
rect 369362 420960 369410 421016
rect 369301 420958 369410 420960
rect 369301 420955 369367 420958
rect 371969 420746 372035 420749
rect 516317 420746 516383 420749
rect 369932 420744 372035 420746
rect 369932 420688 371974 420744
rect 372030 420688 372035 420744
rect 369932 420686 372035 420688
rect 513820 420744 516383 420746
rect 513820 420688 516322 420744
rect 516378 420688 516383 420744
rect 513820 420686 516383 420688
rect 371969 420683 372035 420686
rect 516317 420683 516383 420686
rect 445569 420610 445635 420613
rect 441876 420608 445635 420610
rect 441876 420552 445574 420608
rect 445630 420552 445635 420608
rect 441876 420550 445635 420552
rect 445569 420547 445635 420550
rect 370129 420202 370195 420205
rect 516777 420202 516843 420205
rect 369932 420200 370195 420202
rect 369932 420144 370134 420200
rect 370190 420144 370195 420200
rect 369932 420142 370195 420144
rect 513820 420200 516843 420202
rect 513820 420144 516782 420200
rect 516838 420144 516843 420200
rect 513820 420142 516843 420144
rect 370129 420139 370195 420142
rect 516777 420139 516843 420142
rect 372429 419658 372495 419661
rect 516777 419658 516843 419661
rect 369932 419656 372495 419658
rect 369932 419600 372434 419656
rect 372490 419600 372495 419656
rect 369932 419598 372495 419600
rect 513820 419656 516843 419658
rect 513820 419600 516782 419656
rect 516838 419600 516843 419656
rect 513820 419598 516843 419600
rect 372429 419595 372495 419598
rect 516777 419595 516843 419598
rect 442073 419522 442139 419525
rect 444465 419522 444531 419525
rect 441876 419520 444531 419522
rect 441876 419464 442078 419520
rect 442134 419464 444470 419520
rect 444526 419464 444531 419520
rect 441876 419462 444531 419464
rect 442073 419459 442139 419462
rect 444465 419459 444531 419462
rect 371969 419114 372035 419117
rect 516501 419114 516567 419117
rect 369932 419112 372035 419114
rect 369932 419056 371974 419112
rect 372030 419056 372035 419112
rect 369932 419054 372035 419056
rect 513820 419112 516567 419114
rect 513820 419056 516506 419112
rect 516562 419056 516567 419112
rect 513820 419054 516567 419056
rect 371969 419051 372035 419054
rect 516501 419051 516567 419054
rect 372153 418570 372219 418573
rect 516317 418570 516383 418573
rect 369932 418568 372219 418570
rect 369932 418512 372158 418568
rect 372214 418512 372219 418568
rect 369932 418510 372219 418512
rect 513820 418568 516383 418570
rect 513820 418512 516322 418568
rect 516378 418512 516383 418568
rect 513820 418510 516383 418512
rect 372153 418507 372219 418510
rect 516317 418507 516383 418510
rect 443269 418298 443335 418301
rect 443453 418298 443519 418301
rect 441876 418296 443519 418298
rect 441876 418240 443274 418296
rect 443330 418240 443458 418296
rect 443514 418240 443519 418296
rect 441876 418238 443519 418240
rect 443269 418235 443335 418238
rect 443453 418235 443519 418238
rect 580533 418298 580599 418301
rect 583520 418298 584960 418388
rect 580533 418296 584960 418298
rect 580533 418240 580538 418296
rect 580594 418240 584960 418296
rect 580533 418238 584960 418240
rect 580533 418235 580599 418238
rect 583520 418148 584960 418238
rect 370221 418026 370287 418029
rect 516317 418026 516383 418029
rect 369932 418024 370287 418026
rect 369932 417996 370226 418024
rect 369902 417968 370226 417996
rect 370282 417968 370287 418024
rect 369902 417966 370287 417968
rect 513820 418024 516383 418026
rect 513820 417968 516322 418024
rect 516378 417968 516383 418024
rect 513820 417966 516383 417968
rect 369902 417757 369962 417966
rect 370221 417963 370287 417966
rect 516317 417963 516383 417966
rect 369902 417752 370011 417757
rect 369902 417696 369950 417752
rect 370006 417696 370011 417752
rect 369902 417694 370011 417696
rect 369945 417691 370011 417694
rect 370865 417482 370931 417485
rect 517421 417482 517487 417485
rect 369932 417480 370931 417482
rect 369932 417424 370870 417480
rect 370926 417424 370931 417480
rect 369932 417422 370931 417424
rect 513820 417480 517487 417482
rect 513820 417424 517426 417480
rect 517482 417424 517487 417480
rect 513820 417422 517487 417424
rect 370865 417419 370931 417422
rect 517421 417419 517487 417422
rect 444649 417210 444715 417213
rect 441876 417208 444715 417210
rect 441876 417152 444654 417208
rect 444710 417152 444715 417208
rect 441876 417150 444715 417152
rect 444649 417147 444715 417150
rect 371969 416938 372035 416941
rect 516593 416938 516659 416941
rect 369932 416936 372035 416938
rect 369932 416880 371974 416936
rect 372030 416880 372035 416936
rect 369932 416878 372035 416880
rect 513820 416936 516659 416938
rect 513820 416880 516598 416936
rect 516654 416880 516659 416936
rect 513820 416878 516659 416880
rect 371969 416875 372035 416878
rect 516593 416875 516659 416878
rect 371969 416394 372035 416397
rect 516501 416394 516567 416397
rect 369932 416392 372035 416394
rect 369932 416336 371974 416392
rect 372030 416336 372035 416392
rect 369932 416334 372035 416336
rect 513820 416392 516567 416394
rect 513820 416336 516506 416392
rect 516562 416336 516567 416392
rect 513820 416334 516567 416336
rect 371969 416331 372035 416334
rect 516501 416331 516567 416334
rect 442165 415986 442231 415989
rect 442625 415986 442691 415989
rect 441876 415984 442691 415986
rect 441876 415928 442170 415984
rect 442226 415928 442630 415984
rect 442686 415928 442691 415984
rect 441876 415926 442691 415928
rect 442165 415923 442231 415926
rect 442625 415923 442691 415926
rect 371969 415850 372035 415853
rect 516317 415850 516383 415853
rect 369932 415848 372035 415850
rect 369932 415792 371974 415848
rect 372030 415792 372035 415848
rect 369932 415790 372035 415792
rect 513820 415848 516383 415850
rect 513820 415792 516322 415848
rect 516378 415792 516383 415848
rect 513820 415790 516383 415792
rect 371969 415787 372035 415790
rect 516317 415787 516383 415790
rect 371233 415306 371299 415309
rect 516501 415306 516567 415309
rect 369932 415304 371299 415306
rect 369932 415248 371238 415304
rect 371294 415248 371299 415304
rect 369932 415246 371299 415248
rect 513820 415304 516567 415306
rect 513820 415248 516506 415304
rect 516562 415248 516567 415304
rect 513820 415246 516567 415248
rect 371233 415243 371299 415246
rect 516501 415243 516567 415246
rect 443361 414898 443427 414901
rect 444189 414898 444255 414901
rect 441876 414896 444255 414898
rect 441876 414840 443366 414896
rect 443422 414840 444194 414896
rect 444250 414840 444255 414896
rect 441876 414838 444255 414840
rect 443361 414835 443427 414838
rect 444189 414835 444255 414838
rect 371969 414762 372035 414765
rect 516317 414762 516383 414765
rect 369932 414760 372035 414762
rect 369932 414704 371974 414760
rect 372030 414704 372035 414760
rect 369932 414702 372035 414704
rect 513820 414760 516383 414762
rect 513820 414704 516322 414760
rect 516378 414704 516383 414760
rect 513820 414702 516383 414704
rect 371969 414699 372035 414702
rect 516317 414699 516383 414702
rect 370221 414218 370287 414221
rect 370681 414218 370747 414221
rect 516317 414218 516383 414221
rect 369932 414216 370747 414218
rect 369932 414160 370226 414216
rect 370282 414160 370686 414216
rect 370742 414160 370747 414216
rect 369932 414158 370747 414160
rect 513820 414216 516383 414218
rect 513820 414160 516322 414216
rect 516378 414160 516383 414216
rect 513820 414158 516383 414160
rect 370221 414155 370287 414158
rect 370681 414155 370747 414158
rect 516317 414155 516383 414158
rect 369393 413946 369459 413949
rect 369350 413944 369459 413946
rect 369350 413888 369398 413944
rect 369454 413888 369459 413944
rect 369350 413883 369459 413888
rect 369350 413674 369410 413883
rect 371233 413674 371299 413677
rect 445477 413674 445543 413677
rect 516777 413674 516843 413677
rect 369350 413672 371299 413674
rect 369350 413644 371238 413672
rect 369380 413616 371238 413644
rect 371294 413616 371299 413672
rect 369380 413614 371299 413616
rect 441876 413672 445543 413674
rect 441876 413616 445482 413672
rect 445538 413616 445543 413672
rect 441876 413614 445543 413616
rect 513820 413672 516843 413674
rect 513820 413616 516782 413672
rect 516838 413616 516843 413672
rect 513820 413614 516843 413616
rect 371233 413611 371299 413614
rect 445477 413611 445543 413614
rect 516777 413611 516843 413614
rect 372797 413130 372863 413133
rect 516317 413130 516383 413133
rect 369932 413128 372863 413130
rect 369932 413072 372802 413128
rect 372858 413072 372863 413128
rect 369932 413070 372863 413072
rect 513820 413128 516383 413130
rect 513820 413072 516322 413128
rect 516378 413072 516383 413128
rect 513820 413070 516383 413072
rect 372797 413067 372863 413070
rect 516317 413067 516383 413070
rect 372061 412586 372127 412589
rect 445477 412586 445543 412589
rect 516317 412586 516383 412589
rect 369932 412584 372127 412586
rect 369932 412528 372066 412584
rect 372122 412528 372127 412584
rect 369932 412526 372127 412528
rect 441876 412584 445543 412586
rect 441876 412528 445482 412584
rect 445538 412528 445543 412584
rect 441876 412526 445543 412528
rect 513820 412584 516383 412586
rect 513820 412528 516322 412584
rect 516378 412528 516383 412584
rect 513820 412526 516383 412528
rect 372061 412523 372127 412526
rect 445477 412523 445543 412526
rect 516317 412523 516383 412526
rect 370497 412178 370563 412181
rect 517605 412178 517671 412181
rect 369932 412176 370563 412178
rect 369932 412148 370502 412176
rect 369902 412120 370502 412148
rect 370558 412120 370563 412176
rect 513452 412176 517671 412178
rect 513452 412148 517610 412176
rect 369902 412118 370563 412120
rect 362769 412044 362835 412045
rect 362718 411980 362724 412044
rect 362788 412042 362835 412044
rect 365161 412042 365227 412045
rect 365294 412042 365300 412044
rect 362788 412040 362880 412042
rect 362830 411984 362880 412040
rect 362788 411982 362880 411984
rect 365161 412040 365300 412042
rect 365161 411984 365166 412040
rect 365222 411984 365300 412040
rect 365161 411982 365300 411984
rect 362788 411980 362835 411982
rect 362769 411979 362835 411980
rect 365161 411979 365227 411982
rect 365294 411980 365300 411982
rect 365364 411980 365370 412044
rect 369902 411637 369962 412118
rect 370497 412115 370563 412118
rect 513422 412120 517610 412148
rect 517666 412120 517671 412176
rect 513422 412118 517671 412120
rect 513422 411637 513482 412118
rect 517605 412115 517671 412118
rect 369853 411632 369962 411637
rect 369853 411576 369858 411632
rect 369914 411576 369962 411632
rect 369853 411574 369962 411576
rect 513373 411632 513482 411637
rect 513373 411576 513378 411632
rect 513434 411576 513482 411632
rect 513373 411574 513482 411576
rect 369853 411571 369919 411574
rect 513373 411571 513439 411574
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 440734 409532 440740 409596
rect 440804 409594 440810 409596
rect 441061 409594 441127 409597
rect 440804 409592 441127 409594
rect 440804 409536 441066 409592
rect 441122 409536 441127 409592
rect 440804 409534 441127 409536
rect 440804 409532 440810 409534
rect 441061 409531 441127 409534
rect 361614 409124 361620 409188
rect 361684 409186 361690 409188
rect 362718 409186 362724 409188
rect 361684 409126 362724 409186
rect 361684 409124 361690 409126
rect 362718 409124 362724 409126
rect 362788 409124 362794 409188
rect 434897 408644 434963 408645
rect 434846 408642 434852 408644
rect 434806 408582 434852 408642
rect 434916 408640 434963 408644
rect 434958 408584 434963 408640
rect 434846 408580 434852 408582
rect 434916 408580 434963 408584
rect 436134 408580 436140 408644
rect 436204 408642 436210 408644
rect 436829 408642 436895 408645
rect 436204 408640 436895 408642
rect 436204 408584 436834 408640
rect 436890 408584 436895 408640
rect 436204 408582 436895 408584
rect 436204 408580 436210 408582
rect 434897 408579 434963 408580
rect 436829 408579 436895 408582
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 444925 369746 444991 369749
rect 441692 369744 444991 369746
rect 441692 369716 444930 369744
rect 441662 369688 444930 369716
rect 444986 369688 444991 369744
rect 441662 369686 444991 369688
rect 441662 369477 441722 369686
rect 444925 369683 444991 369686
rect 370957 369474 371023 369477
rect 369932 369472 371023 369474
rect 369932 369416 370962 369472
rect 371018 369416 371023 369472
rect 369932 369414 371023 369416
rect 370957 369411 371023 369414
rect 441613 369472 441722 369477
rect 516133 369474 516199 369477
rect 441613 369416 441618 369472
rect 441674 369416 441722 369472
rect 513820 369472 516199 369474
rect 513820 369444 516138 369472
rect 441613 369414 441722 369416
rect 513790 369416 516138 369444
rect 516194 369416 516199 369472
rect 513790 369414 516199 369416
rect 441613 369411 441679 369414
rect 513790 369205 513850 369414
rect 516133 369411 516199 369414
rect 442257 369202 442323 369205
rect 444833 369202 444899 369205
rect 441876 369200 444899 369202
rect 441876 369144 442262 369200
rect 442318 369144 444838 369200
rect 444894 369144 444899 369200
rect 441876 369142 444899 369144
rect 442257 369139 442323 369142
rect 444833 369139 444899 369142
rect 513741 369200 513850 369205
rect 513741 369144 513746 369200
rect 513802 369144 513850 369200
rect 513741 369142 513850 369144
rect 513741 369139 513807 369142
rect 441337 368930 441403 368933
rect 441294 368928 441403 368930
rect 441294 368872 441342 368928
rect 441398 368872 441403 368928
rect 441294 368867 441403 368872
rect 441294 368658 441354 368867
rect 444373 368658 444439 368661
rect 441294 368656 444439 368658
rect 441294 368628 444378 368656
rect 441324 368600 444378 368628
rect 444434 368600 444439 368656
rect 441324 368598 444439 368600
rect 444373 368595 444439 368598
rect 370589 368386 370655 368389
rect 516133 368386 516199 368389
rect 369932 368384 370655 368386
rect 369932 368328 370594 368384
rect 370650 368328 370655 368384
rect 513820 368384 516199 368386
rect 513820 368356 516138 368384
rect 369932 368326 370655 368328
rect 370589 368323 370655 368326
rect 513790 368328 516138 368356
rect 516194 368328 516199 368384
rect 513790 368326 516199 368328
rect 441294 367845 441354 368084
rect 513649 367978 513715 367981
rect 513790 367978 513850 368326
rect 516133 368323 516199 368326
rect 513649 367976 513850 367978
rect 513649 367920 513654 367976
rect 513710 367920 513850 367976
rect 513649 367918 513850 367920
rect 513649 367915 513715 367918
rect 441294 367840 441403 367845
rect 441294 367784 441342 367840
rect 441398 367784 441403 367840
rect 441294 367782 441403 367784
rect 441337 367779 441403 367782
rect 441613 367842 441679 367845
rect 441613 367840 441906 367842
rect 441613 367784 441618 367840
rect 441674 367784 441906 367840
rect 441613 367782 441906 367784
rect 441613 367779 441679 367782
rect 441846 367570 441906 367782
rect 513741 367706 513807 367709
rect 513741 367704 513850 367706
rect 513741 367648 513746 367704
rect 513802 367648 513850 367704
rect 513741 367643 513850 367648
rect 444598 367570 444604 367572
rect 441846 367540 444604 367570
rect 441876 367510 444604 367540
rect 444598 367508 444604 367510
rect 444668 367508 444674 367572
rect 370313 367162 370379 367165
rect 369932 367160 370379 367162
rect 369932 367104 370318 367160
rect 370374 367104 370379 367160
rect 513790 367162 513850 367643
rect 516133 367162 516199 367165
rect 513790 367160 516199 367162
rect 513790 367132 516138 367160
rect 369932 367102 370379 367104
rect 513820 367104 516138 367132
rect 516194 367104 516199 367160
rect 513820 367102 516199 367104
rect 370313 367099 370379 367102
rect 516133 367099 516199 367102
rect 442257 367026 442323 367029
rect 445385 367026 445451 367029
rect 441876 367024 445451 367026
rect 441876 366968 442262 367024
rect 442318 366968 445390 367024
rect 445446 366968 445451 367024
rect 441876 366966 445451 366968
rect 442257 366963 442323 366966
rect 445385 366963 445451 366966
rect 444281 366482 444347 366485
rect 441876 366480 444347 366482
rect 441876 366424 444286 366480
rect 444342 366424 444347 366480
rect 441876 366422 444347 366424
rect 444281 366419 444347 366422
rect 370957 366074 371023 366077
rect 516409 366074 516475 366077
rect 369932 366072 371023 366074
rect 369932 366016 370962 366072
rect 371018 366016 371023 366072
rect 369932 366014 371023 366016
rect 513820 366072 516475 366074
rect 513820 366016 516414 366072
rect 516470 366016 516475 366072
rect 513820 366014 516475 366016
rect 370957 366011 371023 366014
rect 516409 366011 516475 366014
rect 442441 365938 442507 365941
rect 444649 365938 444715 365941
rect 441876 365936 444715 365938
rect 441876 365880 442446 365936
rect 442502 365880 444654 365936
rect 444710 365880 444715 365936
rect 441876 365878 444715 365880
rect 442441 365875 442507 365878
rect 444649 365875 444715 365878
rect 444189 365394 444255 365397
rect 441876 365392 444255 365394
rect 441876 365336 444194 365392
rect 444250 365336 444255 365392
rect 441876 365334 444255 365336
rect 444189 365331 444255 365334
rect 580625 365122 580691 365125
rect 583520 365122 584960 365212
rect 580625 365120 584960 365122
rect 580625 365064 580630 365120
rect 580686 365064 584960 365120
rect 580625 365062 584960 365064
rect 580625 365059 580691 365062
rect 583520 364972 584960 365062
rect 370957 364850 371023 364853
rect 444925 364850 444991 364853
rect 516225 364850 516291 364853
rect 369932 364848 371023 364850
rect 369932 364792 370962 364848
rect 371018 364792 371023 364848
rect 369932 364790 371023 364792
rect 441876 364848 444991 364850
rect 441876 364792 444930 364848
rect 444986 364792 444991 364848
rect 441876 364790 444991 364792
rect 513820 364848 516291 364850
rect 513820 364792 516230 364848
rect 516286 364792 516291 364848
rect 513820 364790 516291 364792
rect 370957 364787 371023 364790
rect 444925 364787 444991 364790
rect 516225 364787 516291 364790
rect 445569 364306 445635 364309
rect 441876 364304 445635 364306
rect 441876 364248 445574 364304
rect 445630 364248 445635 364304
rect 441876 364246 445635 364248
rect 445569 364243 445635 364246
rect 441705 364034 441771 364037
rect 441662 364032 441771 364034
rect 441662 363976 441710 364032
rect 441766 363976 441771 364032
rect 441662 363971 441771 363976
rect 370405 363762 370471 363765
rect 370773 363762 370839 363765
rect 369932 363760 370839 363762
rect 369932 363704 370410 363760
rect 370466 363704 370778 363760
rect 370834 363704 370839 363760
rect 441662 363732 441722 363971
rect 516133 363762 516199 363765
rect 513820 363760 516199 363762
rect 369932 363702 370839 363704
rect 513820 363704 516138 363760
rect 516194 363704 516199 363760
rect 513820 363702 516199 363704
rect 370405 363699 370471 363702
rect 370773 363699 370839 363702
rect 516133 363699 516199 363702
rect 445109 363218 445175 363221
rect 441876 363216 445175 363218
rect 441876 363160 445114 363216
rect 445170 363160 445175 363216
rect 441876 363158 445175 363160
rect 445109 363155 445175 363158
rect 444465 362674 444531 362677
rect 441876 362672 444531 362674
rect 441876 362616 444470 362672
rect 444526 362616 444531 362672
rect 441876 362614 444531 362616
rect 444465 362611 444531 362614
rect 370957 362538 371023 362541
rect 516133 362538 516199 362541
rect 369932 362536 371023 362538
rect 369932 362480 370962 362536
rect 371018 362480 371023 362536
rect 369932 362478 371023 362480
rect 513820 362536 516199 362538
rect 513820 362480 516138 362536
rect 516194 362480 516199 362536
rect 513820 362478 516199 362480
rect 370957 362475 371023 362478
rect 516133 362475 516199 362478
rect 445109 362130 445175 362133
rect 441876 362128 445175 362130
rect 441876 362072 445114 362128
rect 445170 362072 445175 362128
rect 441876 362070 445175 362072
rect 445109 362067 445175 362070
rect 445109 361586 445175 361589
rect 441876 361584 445175 361586
rect 441876 361528 445114 361584
rect 445170 361528 445175 361584
rect 441876 361526 445175 361528
rect 445109 361523 445175 361526
rect 516777 361450 516843 361453
rect 513820 361448 516843 361450
rect 369902 360906 369962 361420
rect 513820 361392 516782 361448
rect 516838 361392 516843 361448
rect 513820 361390 516843 361392
rect 516777 361387 516843 361390
rect 441613 361314 441679 361317
rect 441613 361312 441722 361314
rect 441613 361256 441618 361312
rect 441674 361256 441722 361312
rect 441613 361251 441722 361256
rect 441662 361012 441722 361251
rect 370037 360906 370103 360909
rect 369902 360904 370103 360906
rect 369902 360848 370042 360904
rect 370098 360848 370103 360904
rect 369902 360846 370103 360848
rect 370037 360843 370103 360846
rect 445109 360498 445175 360501
rect 441876 360496 445175 360498
rect 441876 360440 445114 360496
rect 445170 360440 445175 360496
rect 441876 360438 445175 360440
rect 445109 360435 445175 360438
rect 516133 360226 516199 360229
rect 513820 360224 516199 360226
rect 369350 359821 369410 360196
rect 513820 360168 516138 360224
rect 516194 360168 516199 360224
rect 513820 360166 516199 360168
rect 516133 360163 516199 360166
rect 445385 360090 445451 360093
rect 441876 360088 445451 360090
rect 441876 360032 445390 360088
rect 445446 360032 445451 360088
rect 441876 360030 445451 360032
rect 445385 360027 445451 360030
rect 369301 359816 369410 359821
rect 369301 359760 369306 359816
rect 369362 359760 369410 359816
rect 369301 359758 369410 359760
rect 369301 359755 369367 359758
rect 445109 359546 445175 359549
rect 445293 359546 445359 359549
rect 441876 359544 445359 359546
rect 441876 359488 445114 359544
rect 445170 359488 445298 359544
rect 445354 359488 445359 359544
rect 441876 359486 445359 359488
rect 445109 359483 445175 359486
rect 445293 359483 445359 359486
rect 516133 359138 516199 359141
rect 513820 359136 516199 359138
rect 369718 358869 369778 359108
rect 513820 359080 516138 359136
rect 516194 359080 516199 359136
rect 513820 359078 516199 359080
rect 516133 359075 516199 359078
rect 445017 359002 445083 359005
rect 441876 359000 445083 359002
rect 441876 358944 445022 359000
rect 445078 358944 445083 359000
rect 441876 358942 445083 358944
rect 445017 358939 445083 358942
rect 369718 358864 369827 358869
rect 369718 358808 369766 358864
rect 369822 358808 369827 358864
rect 369718 358806 369827 358808
rect 369761 358803 369827 358806
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect 444741 358458 444807 358461
rect 445201 358458 445267 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect 441876 358456 445267 358458
rect 441876 358400 444746 358456
rect 444802 358400 445206 358456
rect 445262 358400 445267 358456
rect 441876 358398 445267 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 444741 358395 444807 358398
rect 445201 358395 445267 358398
rect 370129 357914 370195 357917
rect 370681 357914 370747 357917
rect 445661 357914 445727 357917
rect 516133 357914 516199 357917
rect 369932 357912 370747 357914
rect 369932 357856 370134 357912
rect 370190 357856 370686 357912
rect 370742 357856 370747 357912
rect 369932 357854 370747 357856
rect 441876 357912 445727 357914
rect 441876 357856 445666 357912
rect 445722 357856 445727 357912
rect 441876 357854 445727 357856
rect 513820 357912 516199 357914
rect 513820 357856 516138 357912
rect 516194 357856 516199 357912
rect 513820 357854 516199 357856
rect 370129 357851 370195 357854
rect 370681 357851 370747 357854
rect 445661 357851 445727 357854
rect 516133 357851 516199 357854
rect 445293 357370 445359 357373
rect 441876 357368 445359 357370
rect 441876 357312 445298 357368
rect 445354 357312 445359 357368
rect 441876 357310 445359 357312
rect 445293 357307 445359 357310
rect 444414 357172 444420 357236
rect 444484 357234 444490 357236
rect 445477 357234 445543 357237
rect 444484 357232 445543 357234
rect 444484 357176 445482 357232
rect 445538 357176 445543 357232
rect 444484 357174 445543 357176
rect 444484 357172 444490 357174
rect 445477 357171 445543 357174
rect 370957 356826 371023 356829
rect 444598 356826 444604 356828
rect 369932 356824 371023 356826
rect 369932 356768 370962 356824
rect 371018 356768 371023 356824
rect 369932 356766 371023 356768
rect 441876 356766 444604 356826
rect 370957 356763 371023 356766
rect 444598 356764 444604 356766
rect 444668 356826 444674 356828
rect 445569 356826 445635 356829
rect 516409 356826 516475 356829
rect 444668 356824 445635 356826
rect 444668 356768 445574 356824
rect 445630 356768 445635 356824
rect 444668 356766 445635 356768
rect 513820 356824 516475 356826
rect 513820 356768 516414 356824
rect 516470 356768 516475 356824
rect 513820 356766 516475 356768
rect 444668 356764 444674 356766
rect 445569 356763 445635 356766
rect 516409 356763 516475 356766
rect 444414 356282 444420 356284
rect 441876 356222 444420 356282
rect 444414 356220 444420 356222
rect 444484 356220 444490 356284
rect 445017 355738 445083 355741
rect 441876 355736 445083 355738
rect 441876 355680 445022 355736
rect 445078 355680 445083 355736
rect 441876 355678 445083 355680
rect 445017 355675 445083 355678
rect 370957 355602 371023 355605
rect 516133 355602 516199 355605
rect 369932 355600 371023 355602
rect 369932 355544 370962 355600
rect 371018 355544 371023 355600
rect 369932 355542 371023 355544
rect 513820 355600 516199 355602
rect 513820 355544 516138 355600
rect 516194 355544 516199 355600
rect 513820 355542 516199 355544
rect 370957 355539 371023 355542
rect 516133 355539 516199 355542
rect 441846 354922 441906 355164
rect 441846 354862 444850 354922
rect 444790 354786 444850 354862
rect 444790 354726 445770 354786
rect 444649 354650 444715 354653
rect 444790 354652 444850 354726
rect 441876 354648 444715 354650
rect 441876 354592 444654 354648
rect 444710 354592 444715 354648
rect 441876 354590 444715 354592
rect 444649 354587 444715 354590
rect 444782 354588 444788 354652
rect 444852 354588 444858 354652
rect 445710 354650 445770 354726
rect 467097 354650 467163 354653
rect 445710 354648 467163 354650
rect 445710 354592 467102 354648
rect 467158 354592 467163 354648
rect 445710 354590 467163 354592
rect 467097 354587 467163 354590
rect 370957 354514 371023 354517
rect 516133 354514 516199 354517
rect 369932 354512 371023 354514
rect 369932 354456 370962 354512
rect 371018 354456 371023 354512
rect 369932 354454 371023 354456
rect 513820 354512 516199 354514
rect 513820 354456 516138 354512
rect 516194 354456 516199 354512
rect 513820 354454 516199 354456
rect 370957 354451 371023 354454
rect 516133 354451 516199 354454
rect 445569 354106 445635 354109
rect 441876 354104 445635 354106
rect 441876 354048 445574 354104
rect 445630 354048 445635 354104
rect 441876 354046 445635 354048
rect 445569 354043 445635 354046
rect 369945 353562 370011 353565
rect 445109 353562 445175 353565
rect 369902 353560 370011 353562
rect 369902 353504 369950 353560
rect 370006 353504 370011 353560
rect 369902 353499 370011 353504
rect 441876 353560 445175 353562
rect 441876 353504 445114 353560
rect 445170 353504 445175 353560
rect 441876 353502 445175 353504
rect 445109 353499 445175 353502
rect 369902 353290 369962 353499
rect 370589 353290 370655 353293
rect 517605 353290 517671 353293
rect 369902 353288 370655 353290
rect 369902 353250 370594 353288
rect 369932 353232 370594 353250
rect 370650 353232 370655 353288
rect 369932 353230 370655 353232
rect 513820 353288 517671 353290
rect 513820 353232 517610 353288
rect 517666 353232 517671 353288
rect 513820 353230 517671 353232
rect 370589 353227 370655 353230
rect 517605 353227 517671 353230
rect 445569 353018 445635 353021
rect 441876 353016 445635 353018
rect 441876 352960 445574 353016
rect 445630 352960 445635 353016
rect 441876 352958 445635 352960
rect 445569 352955 445635 352958
rect 445569 352474 445635 352477
rect 441876 352472 445635 352474
rect 441876 352416 445574 352472
rect 445630 352416 445635 352472
rect 441876 352414 445635 352416
rect 445569 352411 445635 352414
rect 370865 352202 370931 352205
rect 517421 352202 517487 352205
rect 369932 352200 370931 352202
rect 369932 352144 370870 352200
rect 370926 352144 370931 352200
rect 369932 352142 370931 352144
rect 513820 352200 517487 352202
rect 513820 352144 517426 352200
rect 517482 352144 517487 352200
rect 513820 352142 517487 352144
rect 370865 352139 370931 352142
rect 517421 352139 517487 352142
rect 445569 351930 445635 351933
rect 441876 351928 445635 351930
rect 441876 351872 445574 351928
rect 445630 351872 445635 351928
rect 441876 351870 445635 351872
rect 445569 351867 445635 351870
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect 444373 351386 444439 351389
rect 441876 351384 444439 351386
rect 441876 351328 444378 351384
rect 444434 351328 444439 351384
rect 441876 351326 444439 351328
rect 444373 351323 444439 351326
rect 441705 351114 441771 351117
rect 441705 351112 441906 351114
rect 441705 351056 441710 351112
rect 441766 351056 441906 351112
rect 441705 351054 441906 351056
rect 441705 351051 441771 351054
rect 370681 350978 370747 350981
rect 369932 350976 370747 350978
rect 369932 350920 370686 350976
rect 370742 350920 370747 350976
rect 369932 350918 370747 350920
rect 370681 350915 370747 350918
rect 441846 350570 441906 351054
rect 516133 350978 516199 350981
rect 513820 350976 516199 350978
rect 513820 350920 516138 350976
rect 516194 350920 516199 350976
rect 513820 350918 516199 350920
rect 516133 350915 516199 350918
rect 443361 350570 443427 350573
rect 441846 350568 443427 350570
rect 441846 350512 443366 350568
rect 443422 350512 443427 350568
rect 441846 350510 443427 350512
rect 443361 350507 443427 350510
rect 445477 350298 445543 350301
rect 441876 350296 445543 350298
rect 441876 350240 445482 350296
rect 445538 350240 445543 350296
rect 441876 350238 445543 350240
rect 445477 350235 445543 350238
rect 370957 349890 371023 349893
rect 442993 349890 443059 349893
rect 443729 349890 443795 349893
rect 516593 349890 516659 349893
rect 369932 349888 371023 349890
rect 369932 349832 370962 349888
rect 371018 349832 371023 349888
rect 369932 349830 371023 349832
rect 441876 349888 443795 349890
rect 441876 349832 442998 349888
rect 443054 349832 443734 349888
rect 443790 349832 443795 349888
rect 441876 349830 443795 349832
rect 513820 349888 516659 349890
rect 513820 349832 516598 349888
rect 516654 349832 516659 349888
rect 513820 349830 516659 349832
rect 370957 349827 371023 349830
rect 442993 349827 443059 349830
rect 443729 349827 443795 349830
rect 516593 349827 516659 349830
rect 445937 349346 446003 349349
rect 441876 349344 446003 349346
rect 441876 349288 445942 349344
rect 445998 349288 446003 349344
rect 441876 349286 446003 349288
rect 445937 349283 446003 349286
rect 443085 348802 443151 348805
rect 441876 348800 443151 348802
rect 441876 348744 443090 348800
rect 443146 348744 443151 348800
rect 441876 348742 443151 348744
rect 443085 348739 443151 348742
rect 370957 348666 371023 348669
rect 516133 348666 516199 348669
rect 369932 348664 371023 348666
rect 369932 348608 370962 348664
rect 371018 348608 371023 348664
rect 369932 348606 371023 348608
rect 513820 348664 516199 348666
rect 513820 348608 516138 348664
rect 516194 348608 516199 348664
rect 513820 348606 516199 348608
rect 370957 348603 371023 348606
rect 516133 348603 516199 348606
rect 441889 348530 441955 348533
rect 441846 348528 441955 348530
rect 441846 348472 441894 348528
rect 441950 348472 441955 348528
rect 441846 348467 441955 348472
rect 441846 348228 441906 348467
rect 444373 347714 444439 347717
rect 441876 347712 444439 347714
rect 441876 347656 444378 347712
rect 444434 347656 444439 347712
rect 441876 347654 444439 347656
rect 444373 347651 444439 347654
rect 370497 347578 370563 347581
rect 516133 347578 516199 347581
rect 369932 347576 370563 347578
rect 369932 347520 370502 347576
rect 370558 347520 370563 347576
rect 369932 347518 370563 347520
rect 513820 347576 516199 347578
rect 513820 347520 516138 347576
rect 516194 347520 516199 347576
rect 513820 347518 516199 347520
rect 370497 347515 370563 347518
rect 516133 347515 516199 347518
rect 445845 347170 445911 347173
rect 441876 347168 445911 347170
rect 441876 347112 445850 347168
rect 445906 347112 445911 347168
rect 441876 347110 445911 347112
rect 445845 347107 445911 347110
rect 445109 346626 445175 346629
rect 441876 346624 445175 346626
rect 441876 346568 445114 346624
rect 445170 346568 445175 346624
rect 441876 346566 445175 346568
rect 445109 346563 445175 346566
rect 370957 346354 371023 346357
rect 516133 346354 516199 346357
rect 369932 346352 371023 346354
rect 369932 346296 370962 346352
rect 371018 346296 371023 346352
rect 369932 346294 371023 346296
rect 513820 346352 516199 346354
rect 513820 346296 516138 346352
rect 516194 346296 516199 346352
rect 513820 346294 516199 346296
rect 370957 346291 371023 346294
rect 516133 346291 516199 346294
rect 443545 346082 443611 346085
rect 445753 346082 445819 346085
rect 441876 346080 445819 346082
rect 441876 346024 443550 346080
rect 443606 346024 445758 346080
rect 445814 346024 445819 346080
rect 441876 346022 445819 346024
rect 443545 346019 443611 346022
rect 445753 346019 445819 346022
rect 441981 345810 442047 345813
rect 441846 345808 442047 345810
rect 441846 345752 441986 345808
rect 442042 345752 442047 345808
rect 441846 345750 442047 345752
rect 441846 345538 441906 345750
rect 441981 345747 442047 345750
rect 445477 345538 445543 345541
rect 441846 345536 445543 345538
rect 441846 345508 445482 345536
rect -960 345402 480 345492
rect 441876 345480 445482 345508
rect 445538 345480 445543 345536
rect 441876 345478 445543 345480
rect 445477 345475 445543 345478
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 370221 345266 370287 345269
rect 516225 345266 516291 345269
rect 369932 345264 370287 345266
rect 369932 345208 370226 345264
rect 370282 345208 370287 345264
rect 369932 345206 370287 345208
rect 513820 345264 516291 345266
rect 513820 345208 516230 345264
rect 516286 345208 516291 345264
rect 513820 345206 516291 345208
rect 370221 345203 370287 345206
rect 516225 345203 516291 345206
rect 444465 344994 444531 344997
rect 441876 344992 444531 344994
rect 441876 344936 444470 344992
rect 444526 344936 444531 344992
rect 441876 344934 444531 344936
rect 444465 344931 444531 344934
rect 443637 344450 443703 344453
rect 441876 344448 443703 344450
rect 441876 344392 443642 344448
rect 443698 344392 443703 344448
rect 441876 344390 443703 344392
rect 443637 344387 443703 344390
rect 370957 344042 371023 344045
rect 516133 344042 516199 344045
rect 369932 344040 371023 344042
rect 369932 343984 370962 344040
rect 371018 343984 371023 344040
rect 369932 343982 371023 343984
rect 513820 344040 516199 344042
rect 513820 343984 516138 344040
rect 516194 343984 516199 344040
rect 513820 343982 516199 343984
rect 370957 343979 371023 343982
rect 516133 343979 516199 343982
rect 444373 343906 444439 343909
rect 441876 343904 444439 343906
rect 441876 343876 444378 343904
rect 441846 343848 444378 343876
rect 444434 343848 444439 343904
rect 441846 343846 444439 343848
rect 441846 343637 441906 343846
rect 444373 343843 444439 343846
rect 441846 343632 441955 343637
rect 441846 343576 441894 343632
rect 441950 343576 441955 343632
rect 441846 343574 441955 343576
rect 441889 343571 441955 343574
rect 442073 343362 442139 343365
rect 441876 343360 442139 343362
rect 441876 343332 442078 343360
rect 441846 343304 442078 343332
rect 442134 343304 442139 343360
rect 441846 343302 442139 343304
rect 441846 343093 441906 343302
rect 442073 343299 442139 343302
rect 441797 343088 441906 343093
rect 441797 343032 441802 343088
rect 441858 343032 441906 343088
rect 441797 343030 441906 343032
rect 441797 343027 441863 343030
rect 370957 342954 371023 342957
rect 514753 342954 514819 342957
rect 369932 342952 371023 342954
rect 369932 342896 370962 342952
rect 371018 342896 371023 342952
rect 369932 342894 371023 342896
rect 513820 342952 514819 342954
rect 513820 342896 514758 342952
rect 514814 342896 514819 342952
rect 513820 342894 514819 342896
rect 370957 342891 371023 342894
rect 514753 342891 514819 342894
rect 442993 342818 443059 342821
rect 443453 342818 443519 342821
rect 441876 342816 443519 342818
rect 441876 342760 442998 342816
rect 443054 342760 443458 342816
rect 443514 342760 443519 342816
rect 441876 342758 443519 342760
rect 442993 342755 443059 342758
rect 443453 342755 443519 342758
rect 445109 342274 445175 342277
rect 441876 342272 445175 342274
rect 441876 342216 445114 342272
rect 445170 342216 445175 342272
rect 441876 342214 445175 342216
rect 445109 342211 445175 342214
rect 372797 341730 372863 341733
rect 516133 341730 516199 341733
rect 369932 341728 372863 341730
rect 369932 341672 372802 341728
rect 372858 341672 372863 341728
rect 513820 341728 516199 341730
rect 369932 341670 372863 341672
rect 372797 341667 372863 341670
rect 441846 341458 441906 341700
rect 513820 341672 516138 341728
rect 516194 341672 516199 341728
rect 513820 341670 516199 341672
rect 516133 341667 516199 341670
rect 442165 341458 442231 341461
rect 443085 341458 443151 341461
rect 441846 341456 443151 341458
rect 441846 341400 442170 341456
rect 442226 341400 443090 341456
rect 443146 341400 443151 341456
rect 441846 341398 443151 341400
rect 442165 341395 442231 341398
rect 443085 341395 443151 341398
rect 441662 340917 441722 341156
rect 369853 340914 369919 340917
rect 369853 340912 369962 340914
rect 369853 340856 369858 340912
rect 369914 340856 369962 340912
rect 369853 340851 369962 340856
rect 441613 340912 441722 340917
rect 441613 340856 441618 340912
rect 441674 340856 441722 340912
rect 441613 340854 441722 340856
rect 513373 340914 513439 340917
rect 513373 340912 513482 340914
rect 513373 340856 513378 340912
rect 513434 340856 513482 340912
rect 441613 340851 441679 340854
rect 513373 340851 513482 340856
rect 369902 340642 369962 340851
rect 370221 340642 370287 340645
rect 445477 340642 445543 340645
rect 369902 340640 370287 340642
rect 369902 340612 370226 340640
rect 369932 340584 370226 340612
rect 370282 340584 370287 340640
rect 369932 340582 370287 340584
rect 441876 340640 445543 340642
rect 441876 340584 445482 340640
rect 445538 340584 445543 340640
rect 513422 340612 513482 340851
rect 441876 340582 445543 340584
rect 370221 340579 370287 340582
rect 445477 340579 445543 340582
rect 361614 340444 361620 340508
rect 361684 340506 361690 340508
rect 362493 340506 362559 340509
rect 361684 340504 362559 340506
rect 361684 340448 362498 340504
rect 362554 340448 362559 340504
rect 361684 340446 362559 340448
rect 361684 340444 361690 340446
rect 362493 340443 362559 340446
rect 364374 340444 364380 340508
rect 364444 340506 364450 340508
rect 365161 340506 365227 340509
rect 366582 340506 366588 340508
rect 364444 340504 366588 340506
rect 364444 340448 365166 340504
rect 365222 340448 366588 340504
rect 364444 340446 366588 340448
rect 364444 340444 364450 340446
rect 365161 340443 365227 340446
rect 366582 340444 366588 340446
rect 366652 340444 366658 340508
rect 444557 340234 444623 340237
rect 441876 340232 444623 340234
rect 441876 340176 444562 340232
rect 444618 340176 444623 340232
rect 441876 340174 444623 340176
rect 444557 340171 444623 340174
rect 436134 340036 436140 340100
rect 436204 340098 436210 340100
rect 436553 340098 436619 340101
rect 440785 340100 440851 340101
rect 436204 340096 436619 340098
rect 436204 340040 436558 340096
rect 436614 340040 436619 340096
rect 436204 340038 436619 340040
rect 436204 340036 436210 340038
rect 436553 340035 436619 340038
rect 440734 340036 440740 340100
rect 440804 340098 440851 340100
rect 440804 340096 440896 340098
rect 440846 340040 440896 340096
rect 440804 340038 440896 340040
rect 440804 340036 440851 340038
rect 440785 340035 440851 340036
rect 434851 339964 434917 339965
rect 434846 339962 434852 339964
rect 434760 339902 434852 339962
rect 434846 339900 434852 339902
rect 434916 339900 434922 339964
rect 434851 339899 434917 339900
rect 583520 338452 584960 338692
rect 431861 338058 431927 338061
rect 436553 338058 436619 338061
rect 431861 338056 436619 338058
rect 431861 338000 431866 338056
rect 431922 338000 436558 338056
rect 436614 338000 436619 338056
rect 431861 337998 436619 338000
rect 431861 337995 431927 337998
rect 436553 337995 436619 337998
rect 431769 337922 431835 337925
rect 434805 337922 434871 337925
rect 431769 337920 434871 337922
rect 431769 337864 431774 337920
rect 431830 337864 434810 337920
rect 434866 337864 434871 337920
rect 431769 337862 434871 337864
rect 431769 337859 431835 337862
rect 434805 337859 434871 337862
rect -960 332196 480 332436
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 213821 299434 213887 299437
rect 216029 299434 216095 299437
rect 213821 299432 216095 299434
rect 213821 299376 213826 299432
rect 213882 299376 216034 299432
rect 216090 299376 216095 299432
rect 213821 299374 216095 299376
rect 213821 299371 213887 299374
rect 216029 299371 216095 299374
rect 216806 299372 216812 299436
rect 216876 299434 216882 299436
rect 216949 299434 217015 299437
rect 216876 299432 217015 299434
rect 216876 299376 216954 299432
rect 217010 299376 217015 299432
rect 216876 299374 217015 299376
rect 216876 299372 216882 299374
rect 216949 299371 217015 299374
rect 214373 299298 214439 299301
rect 214557 299298 214623 299301
rect 224401 299298 224467 299301
rect 214373 299296 214482 299298
rect 214373 299240 214378 299296
rect 214434 299240 214482 299296
rect 214373 299235 214482 299240
rect 214557 299296 224467 299298
rect 214557 299240 214562 299296
rect 214618 299240 224406 299296
rect 224462 299240 224467 299296
rect 214557 299238 224467 299240
rect 214557 299235 214623 299238
rect 224401 299235 224467 299238
rect 214422 299162 214482 299235
rect 216806 299162 216812 299164
rect 214422 299102 216812 299162
rect 216806 299100 216812 299102
rect 216876 299100 216882 299164
rect 198457 298890 198523 298893
rect 198457 298888 200100 298890
rect 198457 298832 198462 298888
rect 198518 298832 200100 298888
rect 198457 298830 200100 298832
rect 198457 298827 198523 298830
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 302877 298482 302943 298485
rect 299828 298480 302943 298482
rect 299828 298424 302882 298480
rect 302938 298424 302943 298480
rect 299828 298422 302943 298424
rect 302877 298419 302943 298422
rect 400121 298210 400187 298213
rect 516358 298210 516364 298212
rect 400121 298208 516364 298210
rect 400121 298152 400126 298208
rect 400182 298152 516364 298208
rect 400121 298150 516364 298152
rect 400121 298147 400187 298150
rect 516358 298148 516364 298150
rect 516428 298148 516434 298212
rect 371233 298074 371299 298077
rect 371366 298074 371372 298076
rect 371233 298072 371372 298074
rect 371233 298016 371238 298072
rect 371294 298016 371372 298072
rect 371233 298014 371372 298016
rect 371233 298011 371299 298014
rect 371366 298012 371372 298014
rect 371436 298012 371442 298076
rect 371918 298012 371924 298076
rect 371988 298074 371994 298076
rect 372245 298074 372311 298077
rect 371988 298072 372311 298074
rect 371988 298016 372250 298072
rect 372306 298016 372311 298072
rect 371988 298014 372311 298016
rect 371988 298012 371994 298014
rect 372245 298011 372311 298014
rect 371325 297802 371391 297805
rect 516961 297802 517027 297805
rect 369380 297800 371391 297802
rect 369380 297772 371330 297800
rect 369350 297744 371330 297772
rect 371386 297744 371391 297800
rect 513452 297800 517027 297802
rect 513452 297772 516966 297800
rect 369350 297742 371391 297744
rect 369350 297533 369410 297742
rect 371325 297739 371391 297742
rect 513422 297744 516966 297772
rect 517022 297744 517027 297800
rect 513422 297742 517027 297744
rect 513422 297533 513482 297742
rect 516961 297739 517027 297742
rect 369350 297528 369459 297533
rect 444373 297530 444439 297533
rect 369350 297472 369398 297528
rect 369454 297472 369459 297528
rect 441876 297528 444439 297530
rect 441876 297500 444378 297528
rect 369350 297470 369459 297472
rect 369393 297467 369459 297470
rect 441846 297472 444378 297500
rect 444434 297472 444439 297528
rect 441846 297470 444439 297472
rect 369853 297394 369919 297397
rect 369853 297392 369962 297394
rect 369853 297336 369858 297392
rect 369914 297336 369962 297392
rect 369853 297331 369962 297336
rect 369902 297258 369962 297331
rect 371785 297258 371851 297261
rect 369902 297256 371851 297258
rect 369902 297228 371790 297256
rect 369932 297200 371790 297228
rect 371846 297200 371851 297256
rect 369932 297198 371851 297200
rect 371785 297195 371851 297198
rect 441705 296986 441771 296989
rect 441846 296986 441906 297470
rect 444373 297467 444439 297470
rect 513373 297528 513482 297533
rect 513373 297472 513378 297528
rect 513434 297472 513482 297528
rect 513373 297470 513482 297472
rect 513373 297467 513439 297470
rect 517329 297258 517395 297261
rect 513452 297256 517395 297258
rect 513452 297228 517334 297256
rect 441705 296984 441906 296986
rect 441705 296928 441710 296984
rect 441766 296928 441906 296984
rect 441705 296926 441906 296928
rect 513422 297200 517334 297228
rect 517390 297200 517395 297256
rect 513422 297198 517395 297200
rect 441705 296923 441771 296926
rect 513422 296853 513482 297198
rect 517329 297195 517395 297198
rect 198549 296850 198615 296853
rect 198549 296848 200100 296850
rect 198549 296792 198554 296848
rect 198610 296792 200100 296848
rect 198549 296790 200100 296792
rect 513373 296848 513482 296853
rect 513373 296792 513378 296848
rect 513434 296792 513482 296848
rect 513373 296790 513482 296792
rect 198549 296787 198615 296790
rect 513373 296787 513439 296790
rect 371417 296714 371483 296717
rect 517053 296714 517119 296717
rect 369932 296712 371483 296714
rect 369932 296656 371422 296712
rect 371478 296656 371483 296712
rect 513636 296712 517119 296714
rect 513636 296684 517058 296712
rect 369932 296654 371483 296656
rect 371417 296651 371483 296654
rect 513606 296656 517058 296684
rect 517114 296656 517119 296712
rect 513606 296654 517119 296656
rect 444373 296442 444439 296445
rect 441876 296440 444439 296442
rect 441876 296412 444378 296440
rect 441846 296384 444378 296412
rect 444434 296384 444439 296440
rect 441846 296382 444439 296384
rect 372337 296170 372403 296173
rect 372470 296170 372476 296172
rect 369932 296168 372476 296170
rect 369932 296140 372342 296168
rect 369902 296112 372342 296140
rect 372398 296112 372476 296168
rect 369902 296110 372476 296112
rect 369902 295901 369962 296110
rect 372337 296107 372403 296110
rect 372470 296108 372476 296110
rect 372540 296108 372546 296172
rect 441705 296034 441771 296037
rect 441846 296034 441906 296382
rect 444373 296379 444439 296382
rect 513373 296442 513439 296445
rect 513373 296440 513482 296442
rect 513373 296384 513378 296440
rect 513434 296384 513482 296440
rect 513373 296379 513482 296384
rect 513422 296140 513482 296379
rect 513606 296309 513666 296654
rect 517053 296651 517119 296654
rect 513557 296304 513666 296309
rect 513557 296248 513562 296304
rect 513618 296248 513666 296304
rect 513557 296246 513666 296248
rect 513557 296243 513623 296246
rect 441705 296032 441906 296034
rect 441705 295976 441710 296032
rect 441766 295976 441906 296032
rect 441705 295974 441906 295976
rect 441705 295971 441771 295974
rect 369393 295898 369459 295901
rect 369350 295896 369459 295898
rect 369350 295840 369398 295896
rect 369454 295840 369459 295896
rect 369350 295835 369459 295840
rect 369853 295896 369962 295901
rect 513465 295898 513531 295901
rect 516174 295898 516180 295900
rect 369853 295840 369858 295896
rect 369914 295840 369962 295896
rect 369853 295838 369962 295840
rect 513422 295896 516180 295898
rect 513422 295840 513470 295896
rect 513526 295840 516180 295896
rect 513422 295838 516180 295840
rect 369853 295835 369919 295838
rect 513422 295835 513531 295838
rect 516174 295836 516180 295838
rect 516244 295836 516250 295900
rect 369350 295596 369410 295835
rect 513422 295596 513482 295835
rect 302785 295354 302851 295357
rect 299828 295352 302851 295354
rect 299828 295296 302790 295352
rect 302846 295296 302851 295352
rect 299828 295294 302851 295296
rect 302785 295291 302851 295294
rect 371417 295354 371483 295357
rect 371550 295354 371556 295356
rect 371417 295352 371556 295354
rect 371417 295296 371422 295352
rect 371478 295296 371556 295352
rect 371417 295294 371556 295296
rect 371417 295291 371483 295294
rect 371550 295292 371556 295294
rect 371620 295292 371626 295356
rect 371734 295292 371740 295356
rect 371804 295354 371810 295356
rect 372061 295354 372127 295357
rect 371804 295352 372127 295354
rect 371804 295296 372066 295352
rect 372122 295296 372127 295352
rect 371804 295294 372127 295296
rect 371804 295292 371810 295294
rect 372061 295291 372127 295294
rect 445385 295218 445451 295221
rect 441876 295216 445451 295218
rect 441876 295160 445390 295216
rect 445446 295160 445451 295216
rect 441876 295158 445451 295160
rect 445385 295155 445451 295158
rect 370497 295082 370563 295085
rect 371182 295082 371188 295084
rect 369932 295080 371188 295082
rect 369932 295024 370502 295080
rect 370558 295024 371188 295080
rect 369932 295022 371188 295024
rect 370497 295019 370563 295022
rect 371182 295020 371188 295022
rect 371252 295082 371258 295084
rect 372153 295082 372219 295085
rect 516133 295082 516199 295085
rect 371252 295080 372219 295082
rect 371252 295024 372158 295080
rect 372214 295024 372219 295080
rect 371252 295022 372219 295024
rect 513820 295080 516199 295082
rect 513820 295024 516138 295080
rect 516194 295024 516199 295080
rect 513820 295022 516199 295024
rect 371252 295020 371258 295022
rect 372153 295019 372219 295022
rect 516133 295019 516199 295022
rect 198457 294674 198523 294677
rect 198457 294672 200100 294674
rect 198457 294616 198462 294672
rect 198518 294616 200100 294672
rect 198457 294614 200100 294616
rect 198457 294611 198523 294614
rect 370589 294538 370655 294541
rect 371325 294538 371391 294541
rect 516225 294538 516291 294541
rect 369932 294536 371391 294538
rect 369932 294480 370594 294536
rect 370650 294480 371330 294536
rect 371386 294480 371391 294536
rect 369932 294478 371391 294480
rect 513820 294536 516291 294538
rect 513820 294480 516230 294536
rect 516286 294480 516291 294536
rect 513820 294478 516291 294480
rect 370589 294475 370655 294478
rect 371325 294475 371391 294478
rect 516225 294475 516291 294478
rect 445477 294130 445543 294133
rect 441876 294128 445543 294130
rect 441876 294072 445482 294128
rect 445538 294072 445543 294128
rect 441876 294070 445543 294072
rect 445477 294067 445543 294070
rect 371693 293994 371759 293997
rect 516317 293994 516383 293997
rect 369932 293992 371759 293994
rect 369932 293936 371698 293992
rect 371754 293936 371759 293992
rect 369932 293934 371759 293936
rect 513820 293992 516383 293994
rect 513820 293936 516322 293992
rect 516378 293936 516383 293992
rect 513820 293934 516383 293936
rect 371693 293931 371759 293934
rect 516317 293931 516383 293934
rect 516225 293858 516291 293861
rect 516358 293858 516364 293860
rect 516225 293856 516364 293858
rect 516225 293800 516230 293856
rect 516286 293800 516364 293856
rect 516225 293798 516364 293800
rect 516225 293795 516291 293798
rect 516358 293796 516364 293798
rect 516428 293796 516434 293860
rect 371325 293450 371391 293453
rect 516133 293450 516199 293453
rect 369932 293448 371391 293450
rect 369932 293392 371330 293448
rect 371386 293392 371391 293448
rect 369932 293390 371391 293392
rect 513820 293448 516199 293450
rect 513820 293392 516138 293448
rect 516194 293392 516199 293448
rect 513820 293390 516199 293392
rect 371325 293387 371391 293390
rect 516133 293387 516199 293390
rect -960 293178 480 293268
rect 3877 293178 3943 293181
rect -960 293176 3943 293178
rect -960 293120 3882 293176
rect 3938 293120 3943 293176
rect -960 293118 3943 293120
rect -960 293028 480 293118
rect 3877 293115 3943 293118
rect 370681 292906 370747 292909
rect 371233 292906 371299 292909
rect 443637 292906 443703 292909
rect 516225 292906 516291 292909
rect 369932 292904 371299 292906
rect 369932 292848 370686 292904
rect 370742 292848 371238 292904
rect 371294 292848 371299 292904
rect 369932 292846 371299 292848
rect 441876 292904 443703 292906
rect 441876 292848 443642 292904
rect 443698 292848 443703 292904
rect 441876 292846 443703 292848
rect 513820 292904 516291 292906
rect 513820 292848 516230 292904
rect 516286 292848 516291 292904
rect 513820 292846 516291 292848
rect 370681 292843 370747 292846
rect 371233 292843 371299 292846
rect 443637 292843 443703 292846
rect 516225 292843 516291 292846
rect 198641 292634 198707 292637
rect 198641 292632 200100 292634
rect 198641 292576 198646 292632
rect 198702 292576 200100 292632
rect 198641 292574 200100 292576
rect 198641 292571 198707 292574
rect 302969 292362 303035 292365
rect 371233 292362 371299 292365
rect 516133 292362 516199 292365
rect 299828 292360 303035 292362
rect 299828 292304 302974 292360
rect 303030 292304 303035 292360
rect 369932 292360 371299 292362
rect 369932 292332 371238 292360
rect 299828 292302 303035 292304
rect 302969 292299 303035 292302
rect 369902 292304 371238 292332
rect 371294 292304 371299 292360
rect 369902 292302 371299 292304
rect 513820 292360 516199 292362
rect 513820 292304 516138 292360
rect 516194 292304 516199 292360
rect 513820 292302 516199 292304
rect 369485 291954 369551 291957
rect 369902 291954 369962 292302
rect 371233 292299 371299 292302
rect 516133 292299 516199 292302
rect 369485 291952 369962 291954
rect 369485 291896 369490 291952
rect 369546 291896 369962 291952
rect 369485 291894 369962 291896
rect 369485 291891 369551 291894
rect 371693 291818 371759 291821
rect 443361 291818 443427 291821
rect 446489 291818 446555 291821
rect 516317 291818 516383 291821
rect 369932 291816 371759 291818
rect 369932 291760 371698 291816
rect 371754 291760 371759 291816
rect 369932 291758 371759 291760
rect 441876 291816 446555 291818
rect 441876 291760 443366 291816
rect 443422 291760 446494 291816
rect 446550 291760 446555 291816
rect 441876 291758 446555 291760
rect 513820 291816 516383 291818
rect 513820 291760 516322 291816
rect 516378 291760 516383 291816
rect 513820 291758 516383 291760
rect 371693 291755 371759 291758
rect 443361 291755 443427 291758
rect 446489 291755 446555 291758
rect 516317 291755 516383 291758
rect 371693 291274 371759 291277
rect 516225 291274 516291 291277
rect 369932 291272 371759 291274
rect 369932 291216 371698 291272
rect 371754 291216 371759 291272
rect 369932 291214 371759 291216
rect 513820 291272 516291 291274
rect 513820 291216 516230 291272
rect 516286 291216 516291 291272
rect 513820 291214 516291 291216
rect 371693 291211 371759 291214
rect 516225 291211 516291 291214
rect 371693 290730 371759 290733
rect 516225 290730 516291 290733
rect 369932 290728 371759 290730
rect 369932 290672 371698 290728
rect 371754 290672 371759 290728
rect 369932 290670 371759 290672
rect 513820 290728 516291 290730
rect 513820 290672 516230 290728
rect 516286 290672 516291 290728
rect 513820 290670 516291 290672
rect 371693 290667 371759 290670
rect 516225 290667 516291 290670
rect 445477 290594 445543 290597
rect 441876 290592 445543 290594
rect 441876 290536 445482 290592
rect 445538 290536 445543 290592
rect 441876 290534 445543 290536
rect 445477 290531 445543 290534
rect 197353 290458 197419 290461
rect 197353 290456 200100 290458
rect 197353 290400 197358 290456
rect 197414 290400 200100 290456
rect 197353 290398 200100 290400
rect 197353 290395 197419 290398
rect 371785 290186 371851 290189
rect 516317 290186 516383 290189
rect 369932 290184 371851 290186
rect 369932 290128 371790 290184
rect 371846 290128 371851 290184
rect 369932 290126 371851 290128
rect 513820 290184 516383 290186
rect 513820 290128 516322 290184
rect 516378 290128 516383 290184
rect 513820 290126 516383 290128
rect 371785 290123 371851 290126
rect 516317 290123 516383 290126
rect 372286 289852 372292 289916
rect 372356 289914 372362 289916
rect 375097 289914 375163 289917
rect 372356 289912 375163 289914
rect 372356 289856 375102 289912
rect 375158 289856 375163 289912
rect 372356 289854 375163 289856
rect 372356 289852 372362 289854
rect 375097 289851 375163 289854
rect 371233 289642 371299 289645
rect 516133 289642 516199 289645
rect 369932 289640 371299 289642
rect 369932 289584 371238 289640
rect 371294 289584 371299 289640
rect 369932 289582 371299 289584
rect 513820 289640 516199 289642
rect 513820 289584 516138 289640
rect 516194 289584 516199 289640
rect 513820 289582 516199 289584
rect 371233 289579 371299 289582
rect 516133 289579 516199 289582
rect 372102 289444 372108 289508
rect 372172 289506 372178 289508
rect 375189 289506 375255 289509
rect 443545 289506 443611 289509
rect 444281 289506 444347 289509
rect 372172 289504 375255 289506
rect 372172 289448 375194 289504
rect 375250 289448 375255 289504
rect 372172 289446 375255 289448
rect 441876 289504 444347 289506
rect 441876 289448 443550 289504
rect 443606 289448 444286 289504
rect 444342 289448 444347 289504
rect 441876 289446 444347 289448
rect 372172 289444 372178 289446
rect 375189 289443 375255 289446
rect 443545 289443 443611 289446
rect 444281 289443 444347 289446
rect 302233 289234 302299 289237
rect 299828 289232 302299 289234
rect 299828 289176 302238 289232
rect 302294 289176 302299 289232
rect 299828 289174 302299 289176
rect 302233 289171 302299 289174
rect 371693 289098 371759 289101
rect 516225 289098 516291 289101
rect 369932 289096 371759 289098
rect 369932 289040 371698 289096
rect 371754 289040 371759 289096
rect 369932 289038 371759 289040
rect 513820 289096 516291 289098
rect 513820 289040 516230 289096
rect 516286 289040 516291 289096
rect 513820 289038 516291 289040
rect 371693 289035 371759 289038
rect 516225 289035 516291 289038
rect 371693 288554 371759 288557
rect 516317 288554 516383 288557
rect 369932 288552 371759 288554
rect 369932 288496 371698 288552
rect 371754 288496 371759 288552
rect 369932 288494 371759 288496
rect 513820 288552 516383 288554
rect 513820 288496 516322 288552
rect 516378 288496 516383 288552
rect 513820 288494 516383 288496
rect 371693 288491 371759 288494
rect 516317 288491 516383 288494
rect 198549 288418 198615 288421
rect 198549 288416 200100 288418
rect 198549 288360 198554 288416
rect 198610 288360 200100 288416
rect 198549 288358 200100 288360
rect 198549 288355 198615 288358
rect 445937 288282 446003 288285
rect 513925 288282 513991 288285
rect 441876 288280 446003 288282
rect 441876 288224 445942 288280
rect 445998 288224 446003 288280
rect 441876 288222 446003 288224
rect 445937 288219 446003 288222
rect 513790 288280 513991 288282
rect 513790 288224 513930 288280
rect 513986 288224 513991 288280
rect 513790 288222 513991 288224
rect 371877 288146 371943 288149
rect 369932 288144 371943 288146
rect 369932 288116 371882 288144
rect 369902 288088 371882 288116
rect 371938 288088 371943 288144
rect 513790 288116 513850 288222
rect 513925 288219 513991 288222
rect 369902 288086 371943 288088
rect 369902 287877 369962 288086
rect 371877 288083 371943 288086
rect 369902 287872 370011 287877
rect 513649 287874 513715 287877
rect 369902 287816 369950 287872
rect 370006 287816 370011 287872
rect 369902 287814 370011 287816
rect 369945 287811 370011 287814
rect 513606 287872 513715 287874
rect 513606 287816 513654 287872
rect 513710 287816 513715 287872
rect 513606 287811 513715 287816
rect 371325 287602 371391 287605
rect 369932 287600 371391 287602
rect 369932 287544 371330 287600
rect 371386 287544 371391 287600
rect 513606 287572 513666 287811
rect 369932 287542 371391 287544
rect 371325 287539 371391 287542
rect 443177 287194 443243 287197
rect 441876 287192 443243 287194
rect 441876 287136 443182 287192
rect 443238 287136 443243 287192
rect 441876 287134 443243 287136
rect 443177 287131 443243 287134
rect 371509 287058 371575 287061
rect 369932 287056 371575 287058
rect 369932 287000 371514 287056
rect 371570 287000 371575 287056
rect 369932 286998 371575 287000
rect 371509 286995 371575 286998
rect 513790 286789 513850 287028
rect 513557 286786 513623 286789
rect 513557 286784 513666 286786
rect 513557 286728 513562 286784
rect 513618 286728 513666 286784
rect 513557 286723 513666 286728
rect 513790 286784 513899 286789
rect 513790 286728 513838 286784
rect 513894 286728 513899 286784
rect 513790 286726 513899 286728
rect 513833 286723 513899 286726
rect 371969 286514 372035 286517
rect 441981 286514 442047 286517
rect 369932 286512 372035 286514
rect 369932 286456 371974 286512
rect 372030 286456 372035 286512
rect 369932 286454 372035 286456
rect 371969 286451 372035 286454
rect 441846 286512 442047 286514
rect 441846 286456 441986 286512
rect 442042 286456 442047 286512
rect 513606 286484 513666 286723
rect 441846 286454 442047 286456
rect 198181 286242 198247 286245
rect 198181 286240 200100 286242
rect 198181 286184 198186 286240
rect 198242 286184 200100 286240
rect 198181 286182 200100 286184
rect 198181 286179 198247 286182
rect 302233 286106 302299 286109
rect 299828 286104 302299 286106
rect 299828 286048 302238 286104
rect 302294 286048 302299 286104
rect 299828 286046 302299 286048
rect 302233 286043 302299 286046
rect 371141 285970 371207 285973
rect 369932 285968 371207 285970
rect 369932 285912 371146 285968
rect 371202 285912 371207 285968
rect 441846 285940 441906 286454
rect 441981 286451 442047 286454
rect 513373 286242 513439 286245
rect 513373 286240 513482 286242
rect 513373 286184 513378 286240
rect 513434 286184 513482 286240
rect 513373 286179 513482 286184
rect 513422 285940 513482 286179
rect 369932 285910 371207 285912
rect 371141 285907 371207 285910
rect 370405 285426 370471 285429
rect 372337 285426 372403 285429
rect 516409 285426 516475 285429
rect 369932 285424 372403 285426
rect 369932 285368 370410 285424
rect 370466 285368 372342 285424
rect 372398 285368 372403 285424
rect 369932 285366 372403 285368
rect 513820 285424 516475 285426
rect 513820 285368 516414 285424
rect 516470 285368 516475 285424
rect 513820 285366 516475 285368
rect 370405 285363 370471 285366
rect 372337 285363 372403 285366
rect 516409 285363 516475 285366
rect 583520 285276 584960 285516
rect 372429 284882 372495 284885
rect 444741 284882 444807 284885
rect 516777 284882 516843 284885
rect 369932 284880 372495 284882
rect 369932 284852 372434 284880
rect 369902 284824 372434 284852
rect 372490 284824 372495 284880
rect 369902 284822 372495 284824
rect 441876 284880 444807 284882
rect 441876 284824 444746 284880
rect 444802 284824 444807 284880
rect 441876 284822 444807 284824
rect 513820 284880 516843 284882
rect 513820 284824 516782 284880
rect 516838 284824 516843 284880
rect 513820 284822 516843 284824
rect 369902 284477 369962 284822
rect 372429 284819 372495 284822
rect 444741 284819 444807 284822
rect 516777 284819 516843 284822
rect 369853 284472 369962 284477
rect 369853 284416 369858 284472
rect 369914 284416 369962 284472
rect 369853 284414 369962 284416
rect 369853 284411 369919 284414
rect 372245 284338 372311 284341
rect 516501 284338 516567 284341
rect 369932 284336 372311 284338
rect 369932 284280 372250 284336
rect 372306 284280 372311 284336
rect 369932 284278 372311 284280
rect 513820 284336 516567 284338
rect 513820 284280 516506 284336
rect 516562 284280 516567 284336
rect 513820 284278 516567 284280
rect 372245 284275 372311 284278
rect 516501 284275 516567 284278
rect 197353 284202 197419 284205
rect 197353 284200 200100 284202
rect 197353 284144 197358 284200
rect 197414 284144 200100 284200
rect 197353 284142 200100 284144
rect 197353 284139 197419 284142
rect 369342 283868 369348 283932
rect 369412 283868 369418 283932
rect 369350 283389 369410 283868
rect 516409 283794 516475 283797
rect 513820 283792 516475 283794
rect 513820 283736 516414 283792
rect 516470 283736 516475 283792
rect 513820 283734 516475 283736
rect 516409 283731 516475 283734
rect 445845 283658 445911 283661
rect 441876 283656 445911 283658
rect 441876 283600 445850 283656
rect 445906 283600 445911 283656
rect 441876 283598 445911 283600
rect 445845 283595 445911 283598
rect 369350 283384 369459 283389
rect 369350 283328 369398 283384
rect 369454 283328 369459 283384
rect 369350 283326 369459 283328
rect 369393 283323 369459 283326
rect 371509 283250 371575 283253
rect 516593 283250 516659 283253
rect 369932 283248 371575 283250
rect 369932 283192 371514 283248
rect 371570 283192 371575 283248
rect 369932 283190 371575 283192
rect 513820 283248 516659 283250
rect 513820 283192 516598 283248
rect 516654 283192 516659 283248
rect 513820 283190 516659 283192
rect 371509 283187 371575 283190
rect 516593 283187 516659 283190
rect 302785 283114 302851 283117
rect 299828 283112 302851 283114
rect 299828 283056 302790 283112
rect 302846 283056 302851 283112
rect 299828 283054 302851 283056
rect 302785 283051 302851 283054
rect 371601 282706 371667 282709
rect 516317 282706 516383 282709
rect 369932 282704 371667 282706
rect 369932 282648 371606 282704
rect 371662 282648 371667 282704
rect 369932 282646 371667 282648
rect 513820 282704 516383 282706
rect 513820 282648 516322 282704
rect 516378 282648 516383 282704
rect 513820 282646 516383 282648
rect 371601 282643 371667 282646
rect 516317 282643 516383 282646
rect 444373 282570 444439 282573
rect 441876 282568 444439 282570
rect 441876 282512 444378 282568
rect 444434 282512 444439 282568
rect 441876 282510 444439 282512
rect 444373 282507 444439 282510
rect 371693 282162 371759 282165
rect 517145 282162 517211 282165
rect 369932 282160 371759 282162
rect 369932 282104 371698 282160
rect 371754 282104 371759 282160
rect 369932 282102 371759 282104
rect 513820 282160 517211 282162
rect 513820 282104 517150 282160
rect 517206 282104 517211 282160
rect 513820 282102 517211 282104
rect 371693 282099 371759 282102
rect 517145 282099 517211 282102
rect 197905 282026 197971 282029
rect 197905 282024 200100 282026
rect 197905 281968 197910 282024
rect 197966 281968 200100 282024
rect 197905 281966 200100 281968
rect 197905 281963 197971 281966
rect 371233 281618 371299 281621
rect 371509 281618 371575 281621
rect 516133 281618 516199 281621
rect 369932 281616 371575 281618
rect 369932 281560 371238 281616
rect 371294 281560 371514 281616
rect 371570 281560 371575 281616
rect 369932 281558 371575 281560
rect 513820 281616 516199 281618
rect 513820 281560 516138 281616
rect 516194 281560 516199 281616
rect 513820 281558 516199 281560
rect 371233 281555 371299 281558
rect 371509 281555 371575 281558
rect 516133 281555 516199 281558
rect 444741 281346 444807 281349
rect 441876 281344 444807 281346
rect 441876 281288 444746 281344
rect 444802 281288 444807 281344
rect 441876 281286 444807 281288
rect 444741 281283 444807 281286
rect 371509 281074 371575 281077
rect 516225 281074 516291 281077
rect 369932 281072 371575 281074
rect 369932 281016 371514 281072
rect 371570 281016 371575 281072
rect 369932 281014 371575 281016
rect 513820 281072 516291 281074
rect 513820 281016 516230 281072
rect 516286 281016 516291 281072
rect 513820 281014 516291 281016
rect 371509 281011 371575 281014
rect 516225 281011 516291 281014
rect 369393 280802 369459 280805
rect 369350 280800 369459 280802
rect 369350 280744 369398 280800
rect 369454 280744 369459 280800
rect 369350 280739 369459 280744
rect 369350 280500 369410 280739
rect 516133 280530 516199 280533
rect 513820 280528 516199 280530
rect 513820 280472 516138 280528
rect 516194 280472 516199 280528
rect 513820 280470 516199 280472
rect 516133 280467 516199 280470
rect 445477 280258 445543 280261
rect 441876 280256 445543 280258
rect -960 279972 480 280212
rect 441876 280200 445482 280256
rect 445538 280200 445543 280256
rect 441876 280198 445543 280200
rect 445477 280195 445543 280198
rect 444465 280122 444531 280125
rect 445293 280122 445359 280125
rect 444465 280120 445359 280122
rect 444465 280064 444470 280120
rect 444526 280064 445298 280120
rect 445354 280064 445359 280120
rect 444465 280062 445359 280064
rect 444465 280059 444531 280062
rect 445293 280059 445359 280062
rect 197537 279986 197603 279989
rect 302417 279986 302483 279989
rect 371417 279986 371483 279989
rect 516225 279986 516291 279989
rect 197537 279984 200100 279986
rect 197537 279928 197542 279984
rect 197598 279928 200100 279984
rect 197537 279926 200100 279928
rect 299828 279984 302483 279986
rect 299828 279928 302422 279984
rect 302478 279928 302483 279984
rect 299828 279926 302483 279928
rect 369932 279984 371483 279986
rect 369932 279928 371422 279984
rect 371478 279928 371483 279984
rect 369932 279926 371483 279928
rect 513820 279984 516291 279986
rect 513820 279928 516230 279984
rect 516286 279928 516291 279984
rect 513820 279926 516291 279928
rect 197537 279923 197603 279926
rect 302417 279923 302483 279926
rect 371417 279923 371483 279926
rect 516225 279923 516291 279926
rect 371601 279442 371667 279445
rect 516133 279442 516199 279445
rect 369932 279440 371667 279442
rect 369932 279384 371606 279440
rect 371662 279384 371667 279440
rect 369932 279382 371667 279384
rect 513820 279440 516199 279442
rect 513820 279384 516138 279440
rect 516194 279384 516199 279440
rect 513820 279382 516199 279384
rect 371601 279379 371667 279382
rect 516133 279379 516199 279382
rect 445293 279034 445359 279037
rect 441876 279032 445359 279034
rect 441876 278976 445298 279032
rect 445354 278976 445359 279032
rect 441876 278974 445359 278976
rect 445293 278971 445359 278974
rect 370313 278898 370379 278901
rect 370773 278898 370839 278901
rect 517789 278898 517855 278901
rect 369932 278896 370839 278898
rect 369932 278840 370318 278896
rect 370374 278840 370778 278896
rect 370834 278840 370839 278896
rect 369932 278838 370839 278840
rect 513820 278896 517855 278898
rect 513820 278840 517794 278896
rect 517850 278840 517855 278896
rect 513820 278838 517855 278840
rect 370313 278835 370379 278838
rect 370773 278835 370839 278838
rect 517789 278835 517855 278838
rect 371601 278354 371667 278357
rect 516409 278354 516475 278357
rect 369932 278352 371667 278354
rect 369932 278296 371606 278352
rect 371662 278296 371667 278352
rect 369932 278294 371667 278296
rect 513820 278352 516475 278354
rect 513820 278296 516414 278352
rect 516470 278296 516475 278352
rect 513820 278294 516475 278296
rect 371601 278291 371667 278294
rect 516409 278291 516475 278294
rect 370037 278082 370103 278085
rect 372981 278082 373047 278085
rect 369902 278080 373047 278082
rect 369902 278024 370042 278080
rect 370098 278024 372986 278080
rect 373042 278024 373047 278080
rect 369902 278022 373047 278024
rect 369902 277916 369962 278022
rect 370037 278019 370103 278022
rect 372981 278019 373047 278022
rect 444649 277946 444715 277949
rect 516685 277946 516751 277949
rect 441876 277944 444715 277946
rect 441876 277888 444654 277944
rect 444710 277888 444715 277944
rect 441876 277886 444715 277888
rect 513820 277944 516751 277946
rect 513820 277888 516690 277944
rect 516746 277888 516751 277944
rect 513820 277886 516751 277888
rect 444649 277883 444715 277886
rect 516685 277883 516751 277886
rect 197353 277810 197419 277813
rect 197353 277808 200100 277810
rect 197353 277752 197358 277808
rect 197414 277752 200100 277808
rect 197353 277750 200100 277752
rect 197353 277747 197419 277750
rect 369669 277538 369735 277541
rect 369669 277536 369778 277538
rect 369669 277480 369674 277536
rect 369730 277480 369778 277536
rect 369669 277475 369778 277480
rect 369718 277402 369778 277475
rect 371417 277402 371483 277405
rect 516317 277402 516383 277405
rect 369718 277400 371483 277402
rect 369718 277372 371422 277400
rect 369748 277344 371422 277372
rect 371478 277344 371483 277400
rect 369748 277342 371483 277344
rect 513820 277400 516383 277402
rect 513820 277344 516322 277400
rect 516378 277344 516383 277400
rect 513820 277342 516383 277344
rect 371417 277339 371483 277342
rect 516317 277339 516383 277342
rect 370037 276994 370103 276997
rect 369902 276992 370103 276994
rect 369902 276936 370042 276992
rect 370098 276936 370103 276992
rect 369902 276934 370103 276936
rect 302785 276858 302851 276861
rect 299828 276856 302851 276858
rect 299828 276800 302790 276856
rect 302846 276800 302851 276856
rect 369902 276828 369962 276934
rect 370037 276931 370103 276934
rect 516133 276858 516199 276861
rect 513820 276856 516199 276858
rect 299828 276798 302851 276800
rect 513820 276800 516138 276856
rect 516194 276800 516199 276856
rect 513820 276798 516199 276800
rect 302785 276795 302851 276798
rect 516133 276795 516199 276798
rect 444557 276722 444623 276725
rect 441876 276720 444623 276722
rect 441876 276664 444562 276720
rect 444618 276664 444623 276720
rect 441876 276662 444623 276664
rect 444557 276659 444623 276662
rect 372429 276314 372495 276317
rect 516685 276314 516751 276317
rect 369932 276312 372495 276314
rect 369932 276256 372434 276312
rect 372490 276256 372495 276312
rect 369932 276254 372495 276256
rect 513820 276312 516751 276314
rect 513820 276256 516690 276312
rect 516746 276256 516751 276312
rect 513820 276254 516751 276256
rect 372429 276251 372495 276254
rect 516685 276251 516751 276254
rect 197537 275770 197603 275773
rect 371601 275770 371667 275773
rect 197537 275768 200100 275770
rect 197537 275712 197542 275768
rect 197598 275712 200100 275768
rect 197537 275710 200100 275712
rect 369932 275768 371667 275770
rect 369932 275712 371606 275768
rect 371662 275712 371667 275768
rect 369932 275710 371667 275712
rect 197537 275707 197603 275710
rect 371601 275707 371667 275710
rect 441797 275770 441863 275773
rect 516317 275770 516383 275773
rect 441797 275768 441906 275770
rect 441797 275712 441802 275768
rect 441858 275712 441906 275768
rect 441797 275707 441906 275712
rect 513820 275768 516383 275770
rect 513820 275712 516322 275768
rect 516378 275712 516383 275768
rect 513820 275710 516383 275712
rect 516317 275707 516383 275710
rect 441846 275634 441906 275707
rect 445385 275634 445451 275637
rect 441846 275632 445451 275634
rect 441846 275604 445390 275632
rect 441876 275576 445390 275604
rect 445446 275576 445451 275632
rect 441876 275574 445451 275576
rect 445385 275571 445451 275574
rect 372153 275226 372219 275229
rect 516133 275226 516199 275229
rect 369932 275224 372219 275226
rect 369932 275168 372158 275224
rect 372214 275168 372219 275224
rect 369932 275166 372219 275168
rect 513820 275224 516199 275226
rect 513820 275168 516138 275224
rect 516194 275168 516199 275224
rect 513820 275166 516199 275168
rect 372153 275163 372219 275166
rect 516133 275163 516199 275166
rect 372797 274682 372863 274685
rect 516133 274682 516199 274685
rect 369932 274680 372863 274682
rect 369932 274624 372802 274680
rect 372858 274624 372863 274680
rect 369932 274622 372863 274624
rect 513820 274680 516199 274682
rect 513820 274624 516138 274680
rect 516194 274624 516199 274680
rect 513820 274622 516199 274624
rect 372797 274619 372863 274622
rect 516133 274619 516199 274622
rect 442993 274410 443059 274413
rect 444741 274410 444807 274413
rect 441876 274408 444807 274410
rect 441876 274352 442998 274408
rect 443054 274352 444746 274408
rect 444802 274352 444807 274408
rect 441876 274350 444807 274352
rect 442993 274347 443059 274350
rect 444741 274347 444807 274350
rect 371509 274138 371575 274141
rect 516685 274138 516751 274141
rect 369932 274136 371575 274138
rect 369932 274080 371514 274136
rect 371570 274080 371575 274136
rect 369932 274078 371575 274080
rect 513820 274136 516751 274138
rect 513820 274080 516690 274136
rect 516746 274080 516751 274136
rect 513820 274078 516751 274080
rect 371509 274075 371575 274078
rect 516685 274075 516751 274078
rect 302693 273866 302759 273869
rect 299828 273864 302759 273866
rect 299828 273808 302698 273864
rect 302754 273808 302759 273864
rect 299828 273806 302759 273808
rect 302693 273803 302759 273806
rect 197353 273594 197419 273597
rect 371601 273594 371667 273597
rect 517421 273594 517487 273597
rect 197353 273592 200100 273594
rect 197353 273536 197358 273592
rect 197414 273536 200100 273592
rect 197353 273534 200100 273536
rect 369932 273592 371667 273594
rect 369932 273536 371606 273592
rect 371662 273536 371667 273592
rect 369932 273534 371667 273536
rect 513820 273592 517487 273594
rect 513820 273536 517426 273592
rect 517482 273536 517487 273592
rect 513820 273534 517487 273536
rect 197353 273531 197419 273534
rect 371601 273531 371667 273534
rect 517421 273531 517487 273534
rect 444557 273322 444623 273325
rect 441876 273320 444623 273322
rect 441876 273264 444562 273320
rect 444618 273264 444623 273320
rect 441876 273262 444623 273264
rect 444557 273259 444623 273262
rect 371693 273050 371759 273053
rect 516133 273050 516199 273053
rect 369932 273048 371759 273050
rect 369932 272992 371698 273048
rect 371754 272992 371759 273048
rect 369932 272990 371759 272992
rect 513820 273048 516199 273050
rect 513820 272992 516138 273048
rect 516194 272992 516199 273048
rect 513820 272990 516199 272992
rect 371693 272987 371759 272990
rect 516133 272987 516199 272990
rect 371877 272506 371943 272509
rect 516317 272506 516383 272509
rect 369932 272504 371943 272506
rect 369932 272448 371882 272504
rect 371938 272448 371943 272504
rect 369932 272446 371943 272448
rect 513820 272504 516383 272506
rect 513820 272448 516322 272504
rect 516378 272448 516383 272504
rect 513820 272446 516383 272448
rect 371877 272443 371943 272446
rect 516317 272443 516383 272446
rect 580441 272234 580507 272237
rect 583520 272234 584960 272324
rect 580441 272232 584960 272234
rect 580441 272176 580446 272232
rect 580502 272176 584960 272232
rect 580441 272174 584960 272176
rect 580441 272171 580507 272174
rect 443085 272098 443151 272101
rect 441876 272096 443151 272098
rect 441876 272040 443090 272096
rect 443146 272040 443151 272096
rect 583520 272084 584960 272174
rect 441876 272038 443151 272040
rect 443085 272035 443151 272038
rect 371785 271962 371851 271965
rect 516133 271962 516199 271965
rect 369932 271960 371851 271962
rect 369932 271904 371790 271960
rect 371846 271904 371851 271960
rect 369932 271902 371851 271904
rect 513820 271960 516199 271962
rect 513820 271904 516138 271960
rect 516194 271904 516199 271960
rect 513820 271902 516199 271904
rect 371785 271899 371851 271902
rect 516133 271899 516199 271902
rect 197537 271554 197603 271557
rect 441613 271554 441679 271557
rect 197537 271552 200100 271554
rect 197537 271496 197542 271552
rect 197598 271496 200100 271552
rect 197537 271494 200100 271496
rect 441613 271552 441722 271554
rect 441613 271496 441618 271552
rect 441674 271496 441722 271552
rect 197537 271491 197603 271494
rect 441613 271491 441722 271496
rect 372521 271418 372587 271421
rect 369932 271416 372587 271418
rect 369932 271360 372526 271416
rect 372582 271360 372587 271416
rect 369932 271358 372587 271360
rect 372521 271355 372587 271358
rect 441662 270980 441722 271491
rect 516133 271418 516199 271421
rect 513820 271416 516199 271418
rect 513820 271360 516138 271416
rect 516194 271360 516199 271416
rect 513820 271358 516199 271360
rect 516133 271355 516199 271358
rect 371785 270874 371851 270877
rect 516317 270874 516383 270877
rect 369932 270872 371851 270874
rect 369932 270816 371790 270872
rect 371846 270816 371851 270872
rect 369932 270814 371851 270816
rect 513820 270872 516383 270874
rect 513820 270816 516322 270872
rect 516378 270816 516383 270872
rect 513820 270814 516383 270816
rect 371785 270811 371851 270814
rect 516317 270811 516383 270814
rect 303061 270738 303127 270741
rect 299828 270736 303127 270738
rect 299828 270680 303066 270736
rect 303122 270680 303127 270736
rect 299828 270678 303127 270680
rect 303061 270675 303127 270678
rect 371969 270330 372035 270333
rect 516317 270330 516383 270333
rect 369932 270328 372035 270330
rect 369932 270272 371974 270328
rect 372030 270272 372035 270328
rect 369932 270270 372035 270272
rect 513820 270328 516383 270330
rect 513820 270272 516322 270328
rect 516378 270272 516383 270328
rect 513820 270270 516383 270272
rect 371969 270267 372035 270270
rect 516317 270267 516383 270270
rect 371918 269860 371924 269924
rect 371988 269922 371994 269924
rect 372521 269922 372587 269925
rect 371988 269920 372587 269922
rect 371988 269864 372526 269920
rect 372582 269864 372587 269920
rect 371988 269862 372587 269864
rect 371988 269860 371994 269862
rect 372521 269859 372587 269862
rect 371877 269786 371943 269789
rect 445477 269786 445543 269789
rect 516133 269786 516199 269789
rect 369932 269784 371943 269786
rect 369932 269728 371882 269784
rect 371938 269728 371943 269784
rect 369932 269726 371943 269728
rect 441876 269784 445543 269786
rect 441876 269728 445482 269784
rect 445538 269728 445543 269784
rect 441876 269726 445543 269728
rect 513820 269784 516199 269786
rect 513820 269728 516138 269784
rect 516194 269728 516199 269784
rect 513820 269726 516199 269728
rect 371877 269723 371943 269726
rect 445477 269723 445543 269726
rect 516133 269723 516199 269726
rect 198457 269378 198523 269381
rect 198457 269376 200100 269378
rect 198457 269320 198462 269376
rect 198518 269320 200100 269376
rect 198457 269318 200100 269320
rect 198457 269315 198523 269318
rect 371417 269242 371483 269245
rect 516133 269242 516199 269245
rect 369932 269240 371483 269242
rect 369932 269184 371422 269240
rect 371478 269184 371483 269240
rect 369932 269182 371483 269184
rect 513820 269240 516199 269242
rect 513820 269184 516138 269240
rect 516194 269184 516199 269240
rect 513820 269182 516199 269184
rect 371417 269179 371483 269182
rect 516133 269179 516199 269182
rect 372521 268698 372587 268701
rect 445477 268698 445543 268701
rect 516133 268698 516199 268701
rect 369932 268696 372587 268698
rect 369932 268640 372526 268696
rect 372582 268640 372587 268696
rect 369932 268638 372587 268640
rect 441876 268696 445543 268698
rect 441876 268640 445482 268696
rect 445538 268640 445543 268696
rect 441876 268638 445543 268640
rect 513820 268696 516199 268698
rect 513820 268640 516138 268696
rect 516194 268640 516199 268696
rect 513820 268638 516199 268640
rect 372521 268635 372587 268638
rect 445477 268635 445543 268638
rect 516133 268635 516199 268638
rect 513373 268426 513439 268429
rect 513373 268424 513482 268426
rect 513373 268368 513378 268424
rect 513434 268368 513482 268424
rect 513373 268363 513482 268368
rect 513422 268260 513482 268363
rect 369902 268021 369962 268260
rect 369902 268016 370011 268021
rect 369902 267960 369950 268016
rect 370006 267960 370011 268016
rect 369902 267958 370011 267960
rect 369945 267955 370011 267958
rect 302877 267746 302943 267749
rect 299828 267744 302943 267746
rect 299828 267688 302882 267744
rect 302938 267688 302943 267744
rect 299828 267686 302943 267688
rect 302877 267683 302943 267686
rect 444598 267684 444604 267748
rect 444668 267746 444674 267748
rect 449341 267746 449407 267749
rect 444668 267744 449407 267746
rect 444668 267688 449346 267744
rect 449402 267688 449407 267744
rect 444668 267686 449407 267688
rect 444668 267684 444674 267686
rect 449341 267683 449407 267686
rect 197629 267338 197695 267341
rect 197629 267336 200100 267338
rect -960 267202 480 267292
rect 197629 267280 197634 267336
rect 197690 267280 200100 267336
rect 197629 267278 200100 267280
rect 197629 267275 197695 267278
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 358169 266250 358235 266253
rect 361614 266250 361620 266252
rect 358169 266248 361620 266250
rect 358169 266192 358174 266248
rect 358230 266192 361620 266248
rect 358169 266190 361620 266192
rect 358169 266187 358235 266190
rect 361614 266188 361620 266190
rect 361684 266250 361690 266252
rect 362861 266250 362927 266253
rect 361684 266248 362927 266250
rect 361684 266192 362866 266248
rect 362922 266192 362927 266248
rect 361684 266190 362927 266192
rect 361684 266188 361690 266190
rect 362861 266187 362927 266190
rect 356697 266114 356763 266117
rect 356697 266112 364442 266114
rect 356697 266056 356702 266112
rect 356758 266056 364442 266112
rect 356697 266054 364442 266056
rect 356697 266051 356763 266054
rect 364382 265844 364442 266054
rect 364374 265780 364380 265844
rect 364444 265842 364450 265844
rect 364885 265842 364951 265845
rect 364444 265840 364951 265842
rect 364444 265784 364890 265840
rect 364946 265784 364951 265840
rect 364444 265782 364951 265784
rect 364444 265780 364450 265782
rect 364885 265779 364951 265782
rect 436686 265508 436692 265572
rect 436756 265570 436762 265572
rect 436921 265570 436987 265573
rect 436756 265568 436987 265570
rect 436756 265512 436926 265568
rect 436982 265512 436987 265568
rect 436756 265510 436987 265512
rect 436756 265508 436762 265510
rect 436921 265507 436987 265510
rect 197353 265162 197419 265165
rect 197353 265160 200100 265162
rect 197353 265104 197358 265160
rect 197414 265104 200100 265160
rect 197353 265102 200100 265104
rect 197353 265099 197419 265102
rect 434897 265026 434963 265029
rect 435214 265026 435220 265028
rect 434897 265024 435220 265026
rect 434897 264968 434902 265024
rect 434958 264968 435220 265024
rect 434897 264966 435220 264968
rect 434897 264963 434963 264966
rect 435214 264964 435220 264966
rect 435284 264964 435290 265028
rect 302693 264618 302759 264621
rect 299828 264616 302759 264618
rect 299828 264560 302698 264616
rect 302754 264560 302759 264616
rect 299828 264558 302759 264560
rect 302693 264555 302759 264558
rect 197353 263122 197419 263125
rect 197353 263120 200100 263122
rect 197353 263064 197358 263120
rect 197414 263064 200100 263120
rect 197353 263062 200100 263064
rect 197353 263059 197419 263062
rect 302325 261490 302391 261493
rect 299828 261488 302391 261490
rect 299828 261432 302330 261488
rect 302386 261432 302391 261488
rect 299828 261430 302391 261432
rect 302325 261427 302391 261430
rect 197353 260946 197419 260949
rect 197353 260944 200100 260946
rect 197353 260888 197358 260944
rect 197414 260888 200100 260944
rect 197353 260886 200100 260888
rect 197353 260883 197419 260886
rect 197353 258906 197419 258909
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 197353 258904 200100 258906
rect 197353 258848 197358 258904
rect 197414 258848 200100 258904
rect 197353 258846 200100 258848
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 197353 258843 197419 258846
rect 580349 258843 580415 258846
rect 583520 258756 584960 258846
rect 302601 258498 302667 258501
rect 299828 258496 302667 258498
rect 299828 258440 302606 258496
rect 302662 258440 302667 258496
rect 299828 258438 302667 258440
rect 302601 258435 302667 258438
rect 198365 256730 198431 256733
rect 198365 256728 200100 256730
rect 198365 256672 198370 256728
rect 198426 256672 200100 256728
rect 198365 256670 200100 256672
rect 198365 256667 198431 256670
rect 302785 255370 302851 255373
rect 299828 255368 302851 255370
rect 299828 255312 302790 255368
rect 302846 255312 302851 255368
rect 299828 255310 302851 255312
rect 302785 255307 302851 255310
rect 197997 254690 198063 254693
rect 197997 254688 200100 254690
rect 197997 254632 198002 254688
rect 198058 254632 200100 254688
rect 197997 254630 200100 254632
rect 197997 254627 198063 254630
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 197905 252514 197971 252517
rect 197905 252512 200100 252514
rect 197905 252456 197910 252512
rect 197966 252456 200100 252512
rect 197905 252454 200100 252456
rect 197905 252451 197971 252454
rect 302969 252242 303035 252245
rect 303245 252242 303311 252245
rect 299828 252240 303311 252242
rect 299828 252184 302974 252240
rect 303030 252184 303250 252240
rect 303306 252184 303311 252240
rect 299828 252182 303311 252184
rect 302969 252179 303035 252182
rect 303245 252179 303311 252182
rect 198089 250474 198155 250477
rect 198089 250472 200100 250474
rect 198089 250416 198094 250472
rect 198150 250416 200100 250472
rect 198089 250414 200100 250416
rect 198089 250411 198155 250414
rect 302785 249250 302851 249253
rect 299828 249248 302851 249250
rect 299828 249192 302790 249248
rect 302846 249192 302851 249248
rect 299828 249190 302851 249192
rect 302785 249187 302851 249190
rect 197537 248298 197603 248301
rect 197537 248296 200100 248298
rect 197537 248240 197542 248296
rect 197598 248240 200100 248296
rect 197537 248238 200100 248240
rect 197537 248235 197603 248238
rect 198089 246258 198155 246261
rect 198089 246256 200100 246258
rect 198089 246200 198094 246256
rect 198150 246200 200100 246256
rect 198089 246198 200100 246200
rect 198089 246195 198155 246198
rect 302509 246122 302575 246125
rect 299828 246120 302575 246122
rect 299828 246064 302514 246120
rect 302570 246064 302575 246120
rect 299828 246062 302575 246064
rect 302509 246059 302575 246062
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 197537 244082 197603 244085
rect 197537 244080 200100 244082
rect 197537 244024 197542 244080
rect 197598 244024 200100 244080
rect 197537 244022 200100 244024
rect 197537 244019 197603 244022
rect 303245 243130 303311 243133
rect 299828 243128 303311 243130
rect 299828 243072 303250 243128
rect 303306 243072 303311 243128
rect 299828 243070 303311 243072
rect 303245 243067 303311 243070
rect 198273 242042 198339 242045
rect 198273 242040 200100 242042
rect 198273 241984 198278 242040
rect 198334 241984 200100 242040
rect 198273 241982 200100 241984
rect 198273 241979 198339 241982
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 302877 240002 302943 240005
rect 299828 240000 302943 240002
rect 299828 239944 302882 240000
rect 302938 239944 302943 240000
rect 299828 239942 302943 239944
rect 302877 239939 302943 239942
rect 197537 239866 197603 239869
rect 197537 239864 200100 239866
rect 197537 239808 197542 239864
rect 197598 239808 200100 239864
rect 197537 239806 200100 239808
rect 197537 239803 197603 239806
rect 198457 237826 198523 237829
rect 198457 237824 200100 237826
rect 198457 237768 198462 237824
rect 198518 237768 200100 237824
rect 198457 237766 200100 237768
rect 198457 237763 198523 237766
rect 302785 236874 302851 236877
rect 299828 236872 302851 236874
rect 299828 236816 302790 236872
rect 302846 236816 302851 236872
rect 299828 236814 302851 236816
rect 302785 236811 302851 236814
rect 197537 235650 197603 235653
rect 197537 235648 200100 235650
rect 197537 235592 197542 235648
rect 197598 235592 200100 235648
rect 197537 235590 200100 235592
rect 197537 235587 197603 235590
rect 302693 233882 302759 233885
rect 299828 233880 302759 233882
rect 299828 233824 302698 233880
rect 302754 233824 302759 233880
rect 299828 233822 302759 233824
rect 302693 233819 302759 233822
rect 197353 233610 197419 233613
rect 197353 233608 200100 233610
rect 197353 233552 197358 233608
rect 197414 233552 200100 233608
rect 197353 233550 200100 233552
rect 197353 233547 197419 233550
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect 372286 231780 372292 231844
rect 372356 231842 372362 231844
rect 375097 231842 375163 231845
rect 372356 231840 375163 231842
rect 372356 231784 375102 231840
rect 375158 231784 375163 231840
rect 372356 231782 375163 231784
rect 372356 231780 372362 231782
rect 375097 231779 375163 231782
rect 372102 231644 372108 231708
rect 372172 231706 372178 231708
rect 375189 231706 375255 231709
rect 372172 231704 375255 231706
rect 372172 231648 375194 231704
rect 375250 231648 375255 231704
rect 372172 231646 375255 231648
rect 372172 231644 372178 231646
rect 375189 231643 375255 231646
rect 198733 231570 198799 231573
rect 198733 231568 200100 231570
rect 198733 231512 198738 231568
rect 198794 231512 200100 231568
rect 198733 231510 200100 231512
rect 198733 231507 198799 231510
rect 302785 230754 302851 230757
rect 299828 230752 302851 230754
rect 299828 230696 302790 230752
rect 302846 230696 302851 230752
rect 299828 230694 302851 230696
rect 302785 230691 302851 230694
rect 197353 229394 197419 229397
rect 197353 229392 200100 229394
rect 197353 229336 197358 229392
rect 197414 229336 200100 229392
rect 197353 229334 200100 229336
rect 197353 229331 197419 229334
rect -960 227884 480 228124
rect 302785 227626 302851 227629
rect 299828 227624 302851 227626
rect 299828 227568 302790 227624
rect 302846 227568 302851 227624
rect 299828 227566 302851 227568
rect 302785 227563 302851 227566
rect 197537 227354 197603 227357
rect 197537 227352 200100 227354
rect 197537 227296 197542 227352
rect 197598 227296 200100 227352
rect 197537 227294 200100 227296
rect 197537 227291 197603 227294
rect 441613 226266 441679 226269
rect 441613 226264 441722 226266
rect 441613 226208 441618 226264
rect 441674 226208 441722 226264
rect 441613 226203 441722 226208
rect 365110 225660 365116 225724
rect 365180 225722 365186 225724
rect 366582 225722 366588 225724
rect 365180 225662 366588 225722
rect 365180 225660 365186 225662
rect 366582 225660 366588 225662
rect 366652 225660 366658 225724
rect 367829 225722 367895 225725
rect 371233 225722 371299 225725
rect 367829 225720 371299 225722
rect 367829 225664 367834 225720
rect 367890 225664 371238 225720
rect 371294 225664 371299 225720
rect 441662 225692 441722 226203
rect 367829 225662 371299 225664
rect 367829 225659 367895 225662
rect 369350 225420 369410 225662
rect 371233 225659 371299 225662
rect 441613 225586 441679 225589
rect 441613 225584 441722 225586
rect 441613 225528 441618 225584
rect 441674 225528 441722 225584
rect 441613 225523 441722 225528
rect 197353 225178 197419 225181
rect 197353 225176 200100 225178
rect 197353 225120 197358 225176
rect 197414 225120 200100 225176
rect 441662 225148 441722 225523
rect 516133 225450 516199 225453
rect 513820 225448 516199 225450
rect 513820 225420 516138 225448
rect 513790 225392 516138 225420
rect 516194 225392 516199 225448
rect 513790 225390 516199 225392
rect 197353 225118 200100 225120
rect 197353 225115 197419 225118
rect 513790 225045 513850 225390
rect 516133 225387 516199 225390
rect 513741 225040 513850 225045
rect 513741 224984 513746 225040
rect 513802 224984 513850 225040
rect 513741 224982 513850 224984
rect 513741 224979 513807 224982
rect 441613 224906 441679 224909
rect 441613 224904 441722 224906
rect 441613 224848 441618 224904
rect 441674 224848 441722 224904
rect 441613 224843 441722 224848
rect 302325 224634 302391 224637
rect 299828 224632 302391 224634
rect 299828 224576 302330 224632
rect 302386 224576 302391 224632
rect 441662 224604 441722 224843
rect 299828 224574 302391 224576
rect 302325 224571 302391 224574
rect 441705 224498 441771 224501
rect 441662 224496 441771 224498
rect 441662 224440 441710 224496
rect 441766 224440 441771 224496
rect 441662 224435 441771 224440
rect 369350 224229 369410 224332
rect 369350 224224 369459 224229
rect 369350 224168 369398 224224
rect 369454 224168 369459 224224
rect 369350 224166 369459 224168
rect 369393 224163 369459 224166
rect 441662 224060 441722 224435
rect 516133 224362 516199 224365
rect 513820 224360 516199 224362
rect 513820 224332 516138 224360
rect 513790 224304 516138 224332
rect 516194 224304 516199 224360
rect 513790 224302 516199 224304
rect 513790 223957 513850 224302
rect 516133 224299 516199 224302
rect 513741 223952 513850 223957
rect 513741 223896 513746 223952
rect 513802 223896 513850 223952
rect 513741 223894 513850 223896
rect 513741 223891 513807 223894
rect 369485 223682 369551 223685
rect 369485 223680 369594 223682
rect 369485 223624 369490 223680
rect 369546 223624 369594 223680
rect 369485 223619 369594 223624
rect 197997 223138 198063 223141
rect 369534 223138 369594 223619
rect 442073 223546 442139 223549
rect 444741 223546 444807 223549
rect 441876 223544 444807 223546
rect 441876 223488 442078 223544
rect 442134 223488 444746 223544
rect 444802 223488 444807 223544
rect 441876 223486 444807 223488
rect 442073 223483 442139 223486
rect 444741 223483 444807 223486
rect 441981 223410 442047 223413
rect 441846 223408 442047 223410
rect 441846 223352 441986 223408
rect 442042 223352 442047 223408
rect 441846 223350 442047 223352
rect 372521 223138 372587 223141
rect 197997 223136 200100 223138
rect 197997 223080 198002 223136
rect 198058 223080 200100 223136
rect 369534 223136 372587 223138
rect 369534 223108 372526 223136
rect 197997 223078 200100 223080
rect 369564 223080 372526 223108
rect 372582 223080 372587 223136
rect 369564 223078 372587 223080
rect 197997 223075 198063 223078
rect 372521 223075 372587 223078
rect 441846 223002 441906 223350
rect 441981 223347 442047 223350
rect 516593 223138 516659 223141
rect 513820 223136 516659 223138
rect 513820 223080 516598 223136
rect 516654 223080 516659 223136
rect 513820 223078 516659 223080
rect 516593 223075 516659 223078
rect 445661 223002 445727 223005
rect 441846 223000 445727 223002
rect 441846 222972 445666 223000
rect 441876 222944 445666 222972
rect 445722 222944 445727 223000
rect 441876 222942 445727 222944
rect 445661 222939 445727 222942
rect 442349 222458 442415 222461
rect 445569 222458 445635 222461
rect 441876 222456 445635 222458
rect 441876 222400 442354 222456
rect 442410 222400 445574 222456
rect 445630 222400 445635 222456
rect 441876 222398 445635 222400
rect 442349 222395 442415 222398
rect 445569 222395 445635 222398
rect 371509 222050 371575 222053
rect 516133 222050 516199 222053
rect 369932 222048 371575 222050
rect 369932 221992 371514 222048
rect 371570 221992 371575 222048
rect 513452 222048 516199 222050
rect 513452 222020 516138 222048
rect 369932 221990 371575 221992
rect 371509 221987 371575 221990
rect 513422 221992 516138 222020
rect 516194 221992 516199 222048
rect 513422 221990 516199 221992
rect 513422 221917 513482 221990
rect 516133 221987 516199 221990
rect 442165 221914 442231 221917
rect 444741 221914 444807 221917
rect 441876 221912 444807 221914
rect 441876 221856 442170 221912
rect 442226 221856 444746 221912
rect 444802 221856 444807 221912
rect 441876 221854 444807 221856
rect 442165 221851 442231 221854
rect 444741 221851 444807 221854
rect 513373 221912 513482 221917
rect 513373 221856 513378 221912
rect 513434 221856 513482 221912
rect 513373 221854 513482 221856
rect 513373 221851 513439 221854
rect 302325 221506 302391 221509
rect 299828 221504 302391 221506
rect 299828 221448 302330 221504
rect 302386 221448 302391 221504
rect 299828 221446 302391 221448
rect 302325 221443 302391 221446
rect 442257 221370 442323 221373
rect 445569 221370 445635 221373
rect 441876 221368 445635 221370
rect 441876 221312 442262 221368
rect 442318 221312 445574 221368
rect 445630 221312 445635 221368
rect 441876 221310 445635 221312
rect 442257 221307 442323 221310
rect 445569 221307 445635 221310
rect 197353 220962 197419 220965
rect 197353 220960 200100 220962
rect 197353 220904 197358 220960
rect 197414 220904 200100 220960
rect 197353 220902 200100 220904
rect 197353 220899 197419 220902
rect 372337 220826 372403 220829
rect 374729 220826 374795 220829
rect 443545 220826 443611 220829
rect 445661 220826 445727 220829
rect 516133 220826 516199 220829
rect 369932 220824 374795 220826
rect 369932 220768 372342 220824
rect 372398 220768 374734 220824
rect 374790 220768 374795 220824
rect 369932 220766 374795 220768
rect 441876 220824 445727 220826
rect 441876 220768 443550 220824
rect 443606 220768 445666 220824
rect 445722 220768 445727 220824
rect 441876 220766 445727 220768
rect 513820 220824 516199 220826
rect 513820 220768 516138 220824
rect 516194 220768 516199 220824
rect 513820 220766 516199 220768
rect 372337 220763 372403 220766
rect 374729 220763 374795 220766
rect 443545 220763 443611 220766
rect 445661 220763 445727 220766
rect 516133 220763 516199 220766
rect 441797 220690 441863 220693
rect 441797 220688 441906 220690
rect 441797 220632 441802 220688
rect 441858 220632 441906 220688
rect 441797 220627 441906 220632
rect 441846 220282 441906 220627
rect 444741 220282 444807 220285
rect 441846 220280 444807 220282
rect 441846 220252 444746 220280
rect 441876 220224 444746 220252
rect 444802 220224 444807 220280
rect 441876 220222 444807 220224
rect 444741 220219 444807 220222
rect 370313 219738 370379 219741
rect 443085 219738 443151 219741
rect 445569 219738 445635 219741
rect 516133 219738 516199 219741
rect 369932 219736 370379 219738
rect 369932 219680 370318 219736
rect 370374 219680 370379 219736
rect 369932 219678 370379 219680
rect 441876 219736 445635 219738
rect 441876 219680 443090 219736
rect 443146 219680 445574 219736
rect 445630 219680 445635 219736
rect 441876 219678 445635 219680
rect 513820 219736 516199 219738
rect 513820 219680 516138 219736
rect 516194 219680 516199 219736
rect 513820 219678 516199 219680
rect 370313 219675 370379 219678
rect 443085 219675 443151 219678
rect 445569 219675 445635 219678
rect 516133 219675 516199 219678
rect 443637 219194 443703 219197
rect 441876 219192 443703 219194
rect 441876 219136 443642 219192
rect 443698 219136 443703 219192
rect 441876 219134 443703 219136
rect 443637 219131 443703 219134
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 197537 218922 197603 218925
rect 197537 218920 200100 218922
rect 197537 218864 197542 218920
rect 197598 218864 200100 218920
rect 583520 218908 584960 218998
rect 197537 218862 200100 218864
rect 197537 218859 197603 218862
rect 443361 218650 443427 218653
rect 441876 218648 443427 218650
rect 441876 218592 443366 218648
rect 443422 218592 443427 218648
rect 441876 218590 443427 218592
rect 443361 218587 443427 218590
rect 370313 218514 370379 218517
rect 516133 218514 516199 218517
rect 369932 218512 370379 218514
rect 369932 218456 370318 218512
rect 370374 218456 370379 218512
rect 369932 218454 370379 218456
rect 513820 218512 516199 218514
rect 513820 218456 516138 218512
rect 516194 218456 516199 218512
rect 513820 218454 516199 218456
rect 370313 218451 370379 218454
rect 516133 218451 516199 218454
rect 302417 218378 302483 218381
rect 299828 218376 302483 218378
rect 299828 218320 302422 218376
rect 302478 218320 302483 218376
rect 299828 218318 302483 218320
rect 302417 218315 302483 218318
rect 443453 218106 443519 218109
rect 441876 218104 443519 218106
rect 441876 218048 443458 218104
rect 443514 218048 443519 218104
rect 441876 218046 443519 218048
rect 443453 218043 443519 218046
rect 443269 217562 443335 217565
rect 441876 217560 443335 217562
rect 441876 217504 443274 217560
rect 443330 217504 443335 217560
rect 441876 217502 443335 217504
rect 443269 217499 443335 217502
rect 370957 217426 371023 217429
rect 516409 217426 516475 217429
rect 369932 217424 371023 217426
rect 369932 217368 370962 217424
rect 371018 217368 371023 217424
rect 369932 217366 371023 217368
rect 513820 217424 516475 217426
rect 513820 217368 516414 217424
rect 516470 217368 516475 217424
rect 513820 217366 516475 217368
rect 370957 217363 371023 217366
rect 516409 217363 516475 217366
rect 445937 217018 446003 217021
rect 441876 217016 446003 217018
rect 441876 216960 445942 217016
rect 445998 216960 446003 217016
rect 441876 216958 446003 216960
rect 445937 216955 446003 216958
rect 197353 216746 197419 216749
rect 197353 216744 200100 216746
rect 197353 216688 197358 216744
rect 197414 216688 200100 216744
rect 197353 216686 200100 216688
rect 197353 216683 197419 216686
rect 445845 216474 445911 216477
rect 441876 216472 445911 216474
rect 441876 216416 445850 216472
rect 445906 216416 445911 216472
rect 441876 216414 445911 216416
rect 445845 216411 445911 216414
rect 370957 216202 371023 216205
rect 516133 216202 516199 216205
rect 369932 216200 371023 216202
rect 369932 216144 370962 216200
rect 371018 216144 371023 216200
rect 369932 216142 371023 216144
rect 513820 216200 516199 216202
rect 513820 216144 516138 216200
rect 516194 216144 516199 216200
rect 513820 216142 516199 216144
rect 370957 216139 371023 216142
rect 516133 216139 516199 216142
rect 444465 216066 444531 216069
rect 441876 216064 444531 216066
rect 441876 216008 444470 216064
rect 444526 216008 444531 216064
rect 441876 216006 444531 216008
rect 444465 216003 444531 216006
rect 444373 215522 444439 215525
rect 441876 215520 444439 215522
rect 441876 215464 444378 215520
rect 444434 215464 444439 215520
rect 441876 215462 444439 215464
rect 444373 215459 444439 215462
rect 303061 215386 303127 215389
rect 299828 215384 303127 215386
rect 299828 215328 303066 215384
rect 303122 215328 303127 215384
rect 299828 215326 303127 215328
rect 303061 215323 303127 215326
rect 370129 215114 370195 215117
rect 370681 215114 370747 215117
rect 516501 215114 516567 215117
rect 369932 215112 370747 215114
rect -960 214978 480 215068
rect 369932 215056 370134 215112
rect 370190 215056 370686 215112
rect 370742 215056 370747 215112
rect 369932 215054 370747 215056
rect 513820 215112 516567 215114
rect 513820 215056 516506 215112
rect 516562 215056 516567 215112
rect 513820 215054 516567 215056
rect 370129 215051 370195 215054
rect 370681 215051 370747 215054
rect 516501 215051 516567 215054
rect 3325 214978 3391 214981
rect 444557 214978 444623 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect 441876 214976 444623 214978
rect 441876 214920 444562 214976
rect 444618 214920 444623 214976
rect 441876 214918 444623 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 444557 214915 444623 214918
rect 197353 214706 197419 214709
rect 197353 214704 200100 214706
rect 197353 214648 197358 214704
rect 197414 214648 200100 214704
rect 197353 214646 200100 214648
rect 197353 214643 197419 214646
rect 444649 214434 444715 214437
rect 441876 214432 444715 214434
rect 441876 214376 444654 214432
rect 444710 214376 444715 214432
rect 441876 214374 444715 214376
rect 444649 214371 444715 214374
rect 370957 213890 371023 213893
rect 444833 213890 444899 213893
rect 516225 213890 516291 213893
rect 369932 213888 371023 213890
rect 369932 213832 370962 213888
rect 371018 213832 371023 213888
rect 369932 213830 371023 213832
rect 441876 213888 444899 213890
rect 441876 213832 444838 213888
rect 444894 213832 444899 213888
rect 441876 213830 444899 213832
rect 513820 213888 516291 213890
rect 513820 213832 516230 213888
rect 516286 213832 516291 213888
rect 513820 213830 516291 213832
rect 370957 213827 371023 213830
rect 444833 213827 444899 213830
rect 516225 213827 516291 213830
rect 445109 213346 445175 213349
rect 441876 213344 445175 213346
rect 441876 213288 445114 213344
rect 445170 213288 445175 213344
rect 441876 213286 445175 213288
rect 445109 213283 445175 213286
rect 372797 212802 372863 212805
rect 443361 212802 443427 212805
rect 444598 212802 444604 212804
rect 369932 212800 372863 212802
rect 369932 212744 372802 212800
rect 372858 212744 372863 212800
rect 369932 212742 372863 212744
rect 441876 212800 444604 212802
rect 441876 212744 443366 212800
rect 443422 212744 444604 212800
rect 441876 212742 444604 212744
rect 372797 212739 372863 212742
rect 443361 212739 443427 212742
rect 444598 212740 444604 212742
rect 444668 212740 444674 212804
rect 516133 212802 516199 212805
rect 513820 212800 516199 212802
rect 513820 212744 516138 212800
rect 516194 212744 516199 212800
rect 513820 212742 516199 212744
rect 516133 212739 516199 212742
rect 197353 212530 197419 212533
rect 197353 212528 200100 212530
rect 197353 212472 197358 212528
rect 197414 212472 200100 212528
rect 197353 212470 200100 212472
rect 197353 212467 197419 212470
rect 444782 212332 444788 212396
rect 444852 212394 444858 212396
rect 445109 212394 445175 212397
rect 444852 212392 445175 212394
rect 444852 212336 445114 212392
rect 445170 212336 445175 212392
rect 444852 212334 445175 212336
rect 444852 212332 444858 212334
rect 445109 212331 445175 212334
rect 302877 212258 302943 212261
rect 443269 212258 443335 212261
rect 444414 212258 444420 212260
rect 299828 212256 302943 212258
rect 299828 212200 302882 212256
rect 302938 212200 302943 212256
rect 299828 212198 302943 212200
rect 441876 212256 444420 212258
rect 441876 212200 443274 212256
rect 443330 212200 444420 212256
rect 441876 212198 444420 212200
rect 302877 212195 302943 212198
rect 443269 212195 443335 212198
rect 444414 212196 444420 212198
rect 444484 212258 444490 212260
rect 444741 212258 444807 212261
rect 444484 212256 444807 212258
rect 444484 212200 444746 212256
rect 444802 212200 444807 212256
rect 444484 212198 444807 212200
rect 444484 212196 444490 212198
rect 444741 212195 444807 212198
rect 442257 211714 442323 211717
rect 442717 211714 442783 211717
rect 441876 211712 442783 211714
rect 441876 211656 442262 211712
rect 442318 211656 442722 211712
rect 442778 211656 442783 211712
rect 441876 211654 442783 211656
rect 442257 211651 442323 211654
rect 442717 211651 442783 211654
rect 370957 211578 371023 211581
rect 516133 211578 516199 211581
rect 369932 211576 371023 211578
rect 369932 211520 370962 211576
rect 371018 211520 371023 211576
rect 369932 211518 371023 211520
rect 513820 211576 516199 211578
rect 513820 211520 516138 211576
rect 516194 211520 516199 211576
rect 513820 211518 516199 211520
rect 370957 211515 371023 211518
rect 516133 211515 516199 211518
rect 443453 211170 443519 211173
rect 444782 211170 444788 211172
rect 441876 211168 444788 211170
rect 441876 211112 443458 211168
rect 443514 211112 444788 211168
rect 441876 211110 444788 211112
rect 443453 211107 443519 211110
rect 444782 211108 444788 211110
rect 444852 211108 444858 211172
rect 442165 210626 442231 210629
rect 441876 210624 442231 210626
rect 441876 210568 442170 210624
rect 442226 210568 442231 210624
rect 441876 210566 442231 210568
rect 442165 210563 442231 210566
rect 197353 210490 197419 210493
rect 370957 210490 371023 210493
rect 516409 210490 516475 210493
rect 197353 210488 200100 210490
rect 197353 210432 197358 210488
rect 197414 210432 200100 210488
rect 197353 210430 200100 210432
rect 369932 210488 371023 210490
rect 369932 210432 370962 210488
rect 371018 210432 371023 210488
rect 369932 210430 371023 210432
rect 513820 210488 516475 210490
rect 513820 210432 516414 210488
rect 516470 210432 516475 210488
rect 513820 210430 516475 210432
rect 197353 210427 197419 210430
rect 370957 210427 371023 210430
rect 516409 210427 516475 210430
rect 443177 210082 443243 210085
rect 441876 210080 443243 210082
rect 441876 210024 443182 210080
rect 443238 210024 443243 210080
rect 441876 210022 443243 210024
rect 443177 210019 443243 210022
rect 445109 209538 445175 209541
rect 441876 209536 445175 209538
rect 441876 209480 445114 209536
rect 445170 209480 445175 209536
rect 441876 209478 445175 209480
rect 445109 209475 445175 209478
rect 303061 209266 303127 209269
rect 370957 209266 371023 209269
rect 516133 209266 516199 209269
rect 299828 209264 303127 209266
rect 299828 209208 303066 209264
rect 303122 209208 303127 209264
rect 299828 209206 303127 209208
rect 369932 209264 371023 209266
rect 369932 209208 370962 209264
rect 371018 209208 371023 209264
rect 369932 209206 371023 209208
rect 513820 209264 516199 209266
rect 513820 209208 516138 209264
rect 516194 209208 516199 209264
rect 513820 209206 516199 209208
rect 303061 209203 303127 209206
rect 370957 209203 371023 209206
rect 516133 209203 516199 209206
rect 445661 208994 445727 208997
rect 441876 208992 445727 208994
rect 441876 208936 445666 208992
rect 445722 208936 445727 208992
rect 441876 208934 445727 208936
rect 445661 208931 445727 208934
rect 445109 208450 445175 208453
rect 441876 208448 445175 208450
rect 441876 208392 445114 208448
rect 445170 208392 445175 208448
rect 441876 208390 445175 208392
rect 445109 208387 445175 208390
rect 197353 208314 197419 208317
rect 197353 208312 200100 208314
rect 197353 208256 197358 208312
rect 197414 208256 200100 208312
rect 197353 208254 200100 208256
rect 197353 208251 197419 208254
rect 370957 208178 371023 208181
rect 517421 208178 517487 208181
rect 369932 208176 371023 208178
rect 369932 208120 370962 208176
rect 371018 208120 371023 208176
rect 369932 208118 371023 208120
rect 513820 208176 517487 208178
rect 513820 208120 517426 208176
rect 517482 208120 517487 208176
rect 513820 208118 517487 208120
rect 370957 208115 371023 208118
rect 517421 208115 517487 208118
rect 444741 207906 444807 207909
rect 445661 207906 445727 207909
rect 441876 207904 445727 207906
rect 441876 207848 444746 207904
rect 444802 207848 445666 207904
rect 445722 207848 445727 207904
rect 441876 207846 445727 207848
rect 444741 207843 444807 207846
rect 445661 207843 445727 207846
rect 444281 207362 444347 207365
rect 441876 207360 444347 207362
rect 441876 207304 444286 207360
rect 444342 207304 444347 207360
rect 441876 207302 444347 207304
rect 444281 207299 444347 207302
rect 371785 206954 371851 206957
rect 516133 206954 516199 206957
rect 369932 206952 371851 206954
rect 369932 206896 371790 206952
rect 371846 206896 371851 206952
rect 369932 206894 371851 206896
rect 513820 206952 516199 206954
rect 513820 206896 516138 206952
rect 516194 206896 516199 206952
rect 513820 206894 516199 206896
rect 371785 206891 371851 206894
rect 516133 206891 516199 206894
rect 445109 206818 445175 206821
rect 446857 206818 446923 206821
rect 441876 206816 446923 206818
rect 441876 206760 445114 206816
rect 445170 206760 446862 206816
rect 446918 206760 446923 206816
rect 441876 206758 446923 206760
rect 445109 206755 445175 206758
rect 446857 206755 446923 206758
rect 197353 206274 197419 206277
rect 444189 206274 444255 206277
rect 197353 206272 200100 206274
rect 197353 206216 197358 206272
rect 197414 206216 200100 206272
rect 197353 206214 200100 206216
rect 441876 206272 444255 206274
rect 441876 206216 444194 206272
rect 444250 206216 444255 206272
rect 441876 206214 444255 206216
rect 197353 206211 197419 206214
rect 444189 206211 444255 206214
rect 302233 206138 302299 206141
rect 299828 206136 302299 206138
rect 299828 206080 302238 206136
rect 302294 206080 302299 206136
rect 299828 206078 302299 206080
rect 302233 206075 302299 206078
rect 371233 205866 371299 205869
rect 372245 205866 372311 205869
rect 442073 205866 442139 205869
rect 444373 205866 444439 205869
rect 516133 205866 516199 205869
rect 369932 205864 372311 205866
rect 369932 205808 371238 205864
rect 371294 205808 372250 205864
rect 372306 205808 372311 205864
rect 369932 205806 372311 205808
rect 441876 205864 444439 205866
rect 441876 205808 442078 205864
rect 442134 205808 444378 205864
rect 444434 205808 444439 205864
rect 441876 205806 444439 205808
rect 513820 205864 516199 205866
rect 513820 205808 516138 205864
rect 516194 205808 516199 205864
rect 513820 205806 516199 205808
rect 371233 205803 371299 205806
rect 372245 205803 372311 205806
rect 442073 205803 442139 205806
rect 444373 205803 444439 205806
rect 516133 205803 516199 205806
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 442901 205322 442967 205325
rect 441876 205320 442967 205322
rect 441876 205292 442906 205320
rect 441846 205264 442906 205292
rect 442962 205264 442967 205320
rect 441846 205262 442967 205264
rect 441613 205050 441679 205053
rect 441846 205050 441906 205262
rect 442901 205259 442967 205262
rect 441613 205048 441906 205050
rect 441613 204992 441618 205048
rect 441674 204992 441906 205048
rect 441613 204990 441906 204992
rect 441613 204987 441679 204990
rect 444373 204778 444439 204781
rect 441876 204776 444439 204778
rect 441876 204748 444378 204776
rect 441846 204720 444378 204748
rect 444434 204720 444439 204776
rect 441846 204718 444439 204720
rect 441846 204645 441906 204718
rect 444373 204715 444439 204718
rect 372245 204642 372311 204645
rect 369932 204640 372311 204642
rect 369932 204584 372250 204640
rect 372306 204584 372311 204640
rect 369932 204582 372311 204584
rect 372245 204579 372311 204582
rect 441797 204640 441906 204645
rect 516133 204642 516199 204645
rect 441797 204584 441802 204640
rect 441858 204584 441906 204640
rect 441797 204582 441906 204584
rect 513820 204640 516199 204642
rect 513820 204584 516138 204640
rect 516194 204584 516199 204640
rect 513820 204582 516199 204584
rect 441797 204579 441863 204582
rect 516133 204579 516199 204582
rect 445569 204234 445635 204237
rect 441876 204232 445635 204234
rect 441876 204176 445574 204232
rect 445630 204176 445635 204232
rect 441876 204174 445635 204176
rect 445569 204171 445635 204174
rect 198273 204098 198339 204101
rect 198273 204096 200100 204098
rect 198273 204040 198278 204096
rect 198334 204040 200100 204096
rect 198273 204038 200100 204040
rect 198273 204035 198339 204038
rect 442717 203690 442783 203693
rect 441876 203688 442783 203690
rect 441876 203660 442722 203688
rect 441846 203632 442722 203660
rect 442778 203632 442783 203688
rect 441846 203630 442783 203632
rect 371918 203554 371924 203556
rect 369932 203494 371924 203554
rect 371918 203492 371924 203494
rect 371988 203554 371994 203556
rect 372153 203554 372219 203557
rect 371988 203552 372219 203554
rect 371988 203496 372158 203552
rect 372214 203496 372219 203552
rect 371988 203494 372219 203496
rect 441846 203554 441906 203630
rect 442717 203627 442783 203630
rect 441981 203554 442047 203557
rect 516133 203554 516199 203557
rect 441846 203552 442047 203554
rect 441846 203496 441986 203552
rect 442042 203496 442047 203552
rect 441846 203494 442047 203496
rect 513820 203552 516199 203554
rect 513820 203496 516138 203552
rect 516194 203496 516199 203552
rect 513820 203494 516199 203496
rect 371988 203492 371994 203494
rect 372153 203491 372219 203494
rect 441981 203491 442047 203494
rect 516133 203491 516199 203494
rect 442349 203146 442415 203149
rect 441876 203144 442415 203146
rect 441876 203088 442354 203144
rect 442410 203088 442415 203144
rect 441876 203086 442415 203088
rect 442349 203083 442415 203086
rect 302969 203010 303035 203013
rect 299828 203008 303035 203010
rect 299828 202952 302974 203008
rect 303030 202952 303035 203008
rect 299828 202950 303035 202952
rect 302969 202947 303035 202950
rect 445661 202602 445727 202605
rect 441876 202600 445727 202602
rect 441876 202544 445666 202600
rect 445722 202544 445727 202600
rect 441876 202542 445727 202544
rect 445661 202539 445727 202542
rect 371325 202330 371391 202333
rect 372061 202330 372127 202333
rect 516133 202330 516199 202333
rect 369932 202328 372127 202330
rect 369932 202272 371330 202328
rect 371386 202272 372066 202328
rect 372122 202272 372127 202328
rect 369932 202270 372127 202272
rect 513820 202328 516199 202330
rect 513820 202272 516138 202328
rect 516194 202272 516199 202328
rect 513820 202270 516199 202272
rect 371325 202267 371391 202270
rect 372061 202267 372127 202270
rect 516133 202267 516199 202270
rect 197353 202058 197419 202061
rect 442901 202058 442967 202061
rect 197353 202056 200100 202058
rect -960 201922 480 202012
rect 197353 202000 197358 202056
rect 197414 202000 200100 202056
rect 441876 202056 442967 202058
rect 441876 202028 442906 202056
rect 197353 201998 200100 202000
rect 441846 202000 442906 202028
rect 442962 202000 442967 202056
rect 441846 201998 442967 202000
rect 197353 201995 197419 201998
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 441705 201922 441771 201925
rect 441846 201922 441906 201998
rect 442901 201995 442967 201998
rect 441705 201920 441906 201922
rect 441705 201864 441710 201920
rect 441766 201864 441906 201920
rect 441705 201862 441906 201864
rect 441705 201859 441771 201862
rect 445661 201514 445727 201517
rect 441876 201512 445727 201514
rect 441876 201456 445666 201512
rect 445722 201456 445727 201512
rect 441876 201454 445727 201456
rect 445661 201451 445727 201454
rect 444833 201378 444899 201381
rect 445201 201378 445267 201381
rect 444833 201376 445267 201378
rect 444833 201320 444838 201376
rect 444894 201320 445206 201376
rect 445262 201320 445267 201376
rect 444833 201318 445267 201320
rect 444833 201315 444899 201318
rect 445201 201315 445267 201318
rect 371509 201242 371575 201245
rect 371969 201242 372035 201245
rect 444414 201242 444420 201244
rect 369932 201240 372035 201242
rect 369932 201184 371514 201240
rect 371570 201184 371974 201240
rect 372030 201184 372035 201240
rect 369932 201182 372035 201184
rect 371509 201179 371575 201182
rect 371969 201179 372035 201182
rect 441846 201182 444420 201242
rect 441846 200940 441906 201182
rect 444414 201180 444420 201182
rect 444484 201242 444490 201244
rect 445293 201242 445359 201245
rect 514661 201242 514727 201245
rect 444484 201240 445359 201242
rect 444484 201184 445298 201240
rect 445354 201184 445359 201240
rect 513820 201240 514727 201242
rect 513820 201212 514666 201240
rect 444484 201182 445359 201184
rect 444484 201180 444490 201182
rect 445293 201179 445359 201182
rect 513790 201184 514666 201212
rect 514722 201184 514727 201240
rect 513790 201182 514727 201184
rect 513557 200834 513623 200837
rect 513790 200834 513850 201182
rect 514661 201179 514727 201182
rect 513557 200832 513850 200834
rect 513557 200776 513562 200832
rect 513618 200776 513850 200832
rect 513557 200774 513850 200776
rect 513557 200771 513623 200774
rect 444833 200426 444899 200429
rect 441876 200424 444899 200426
rect 441876 200368 444838 200424
rect 444894 200368 444899 200424
rect 441876 200366 444899 200368
rect 444833 200363 444899 200366
rect 303429 200018 303495 200021
rect 371601 200018 371667 200021
rect 514109 200018 514175 200021
rect 299828 200016 303495 200018
rect 299828 199960 303434 200016
rect 303490 199960 303495 200016
rect 299828 199958 303495 199960
rect 369932 200016 371667 200018
rect 369932 199960 371606 200016
rect 371662 199960 371667 200016
rect 513452 200016 514175 200018
rect 513452 199988 514114 200016
rect 369932 199958 371667 199960
rect 303429 199955 303495 199958
rect 371601 199955 371667 199958
rect 513422 199960 514114 199988
rect 514170 199960 514175 200016
rect 513422 199958 514175 199960
rect 197537 199882 197603 199885
rect 445477 199882 445543 199885
rect 197537 199880 200100 199882
rect 197537 199824 197542 199880
rect 197598 199824 200100 199880
rect 197537 199822 200100 199824
rect 441876 199880 445543 199882
rect 441876 199824 445482 199880
rect 445538 199824 445543 199880
rect 441876 199822 445543 199824
rect 197537 199819 197603 199822
rect 445477 199819 445543 199822
rect 513422 199477 513482 199958
rect 514109 199955 514175 199958
rect 513373 199472 513482 199477
rect 513373 199416 513378 199472
rect 513434 199416 513482 199472
rect 513373 199414 513482 199416
rect 513373 199411 513439 199414
rect 441846 199066 441906 199308
rect 441846 199006 444666 199066
rect 371417 198930 371483 198933
rect 444606 198932 444666 199006
rect 369932 198928 371483 198930
rect 369932 198872 371422 198928
rect 371478 198872 371483 198928
rect 369932 198870 371483 198872
rect 371417 198867 371483 198870
rect 444598 198868 444604 198932
rect 444668 198930 444674 198932
rect 445201 198930 445267 198933
rect 514201 198930 514267 198933
rect 444668 198928 445267 198930
rect 444668 198872 445206 198928
rect 445262 198872 445267 198928
rect 444668 198870 445267 198872
rect 513820 198928 514267 198930
rect 513820 198872 514206 198928
rect 514262 198872 514267 198928
rect 513820 198870 514267 198872
rect 444668 198868 444674 198870
rect 445201 198867 445267 198870
rect 514201 198867 514267 198870
rect 444465 198794 444531 198797
rect 444925 198794 444991 198797
rect 441876 198792 444991 198794
rect 441876 198736 444470 198792
rect 444526 198736 444930 198792
rect 444986 198736 444991 198792
rect 441876 198734 444991 198736
rect 444465 198731 444531 198734
rect 444925 198731 444991 198734
rect 445293 198250 445359 198253
rect 441876 198248 445359 198250
rect 441876 198192 445298 198248
rect 445354 198192 445359 198248
rect 441876 198190 445359 198192
rect 445293 198187 445359 198190
rect 197353 197842 197419 197845
rect 197353 197840 200100 197842
rect 197353 197784 197358 197840
rect 197414 197784 200100 197840
rect 197353 197782 200100 197784
rect 197353 197779 197419 197782
rect 370957 197706 371023 197709
rect 442993 197706 443059 197709
rect 445293 197706 445359 197709
rect 514109 197706 514175 197709
rect 369932 197704 371023 197706
rect 369932 197648 370962 197704
rect 371018 197648 371023 197704
rect 369932 197646 371023 197648
rect 441876 197704 445359 197706
rect 441876 197648 442998 197704
rect 443054 197648 445298 197704
rect 445354 197648 445359 197704
rect 441876 197646 445359 197648
rect 513820 197704 514175 197706
rect 513820 197648 514114 197704
rect 514170 197648 514175 197704
rect 513820 197646 514175 197648
rect 370957 197643 371023 197646
rect 442993 197643 443059 197646
rect 445293 197643 445359 197646
rect 514109 197643 514175 197646
rect 445661 197162 445727 197165
rect 441876 197160 445727 197162
rect 441876 197104 445666 197160
rect 445722 197104 445727 197160
rect 441876 197102 445727 197104
rect 445661 197099 445727 197102
rect 302785 196890 302851 196893
rect 369945 196890 370011 196893
rect 299828 196888 302851 196890
rect 299828 196832 302790 196888
rect 302846 196832 302851 196888
rect 299828 196830 302851 196832
rect 302785 196827 302851 196830
rect 369902 196888 370011 196890
rect 369902 196832 369950 196888
rect 370006 196832 370011 196888
rect 369902 196827 370011 196832
rect 369902 196618 369962 196827
rect 370865 196618 370931 196621
rect 445385 196618 445451 196621
rect 517421 196618 517487 196621
rect 369902 196616 370931 196618
rect 369902 196588 370870 196616
rect 369932 196560 370870 196588
rect 370926 196560 370931 196616
rect 369932 196558 370931 196560
rect 441876 196616 445451 196618
rect 441876 196560 445390 196616
rect 445446 196560 445451 196616
rect 441876 196558 445451 196560
rect 513820 196616 517487 196618
rect 513820 196560 517426 196616
rect 517482 196560 517487 196616
rect 513820 196558 517487 196560
rect 370865 196555 370931 196558
rect 445385 196555 445451 196558
rect 517421 196555 517487 196558
rect 365161 196482 365227 196485
rect 365294 196482 365300 196484
rect 365161 196480 365300 196482
rect 365161 196424 365166 196480
rect 365222 196424 365300 196480
rect 365161 196422 365300 196424
rect 365161 196419 365227 196422
rect 365294 196420 365300 196422
rect 365364 196482 365370 196484
rect 366582 196482 366588 196484
rect 365364 196422 366588 196482
rect 365364 196420 365370 196422
rect 366582 196420 366588 196422
rect 366652 196420 366658 196484
rect 445845 196210 445911 196213
rect 441876 196208 445911 196210
rect 441876 196152 445850 196208
rect 445906 196152 445911 196208
rect 441876 196150 445911 196152
rect 445845 196147 445911 196150
rect 435173 196076 435239 196077
rect 436737 196076 436803 196077
rect 435173 196072 435220 196076
rect 435284 196074 435290 196076
rect 436686 196074 436692 196076
rect 435173 196016 435178 196072
rect 435173 196012 435220 196016
rect 435284 196014 435330 196074
rect 436646 196014 436692 196074
rect 436756 196072 436803 196076
rect 436798 196016 436803 196072
rect 435284 196012 435290 196014
rect 436686 196012 436692 196014
rect 436756 196012 436803 196016
rect 435173 196011 435239 196012
rect 436737 196011 436803 196012
rect 197537 195666 197603 195669
rect 197537 195664 200100 195666
rect 197537 195608 197542 195664
rect 197598 195608 200100 195664
rect 197537 195606 200100 195608
rect 197537 195603 197603 195606
rect 361614 194516 361620 194580
rect 361684 194578 361690 194580
rect 362718 194578 362724 194580
rect 361684 194518 362724 194578
rect 361684 194516 361690 194518
rect 362718 194516 362724 194518
rect 362788 194578 362794 194580
rect 362861 194578 362927 194581
rect 362788 194576 362927 194578
rect 362788 194520 362866 194576
rect 362922 194520 362927 194576
rect 362788 194518 362927 194520
rect 362788 194516 362794 194518
rect 362861 194515 362927 194518
rect 302601 193762 302667 193765
rect 299828 193760 302667 193762
rect 299828 193704 302606 193760
rect 302662 193704 302667 193760
rect 299828 193702 302667 193704
rect 302601 193699 302667 193702
rect 197353 193626 197419 193629
rect 197353 193624 200100 193626
rect 197353 193568 197358 193624
rect 197414 193568 200100 193624
rect 197353 193566 200100 193568
rect 197353 193563 197419 193566
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 198273 191450 198339 191453
rect 198273 191448 200100 191450
rect 198273 191392 198278 191448
rect 198334 191392 200100 191448
rect 198273 191390 200100 191392
rect 198273 191387 198339 191390
rect 302417 190770 302483 190773
rect 299828 190768 302483 190770
rect 299828 190712 302422 190768
rect 302478 190712 302483 190768
rect 299828 190710 302483 190712
rect 302417 190707 302483 190710
rect 172421 189954 172487 189957
rect 169894 189952 172487 189954
rect 169894 189896 172426 189952
rect 172482 189896 172487 189952
rect 169894 189894 172487 189896
rect 169894 189448 169954 189894
rect 172421 189891 172487 189894
rect 197353 189410 197419 189413
rect 197353 189408 200100 189410
rect 197353 189352 197358 189408
rect 197414 189352 200100 189408
rect 197353 189350 200100 189352
rect 197353 189347 197419 189350
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 172421 188730 172487 188733
rect 169894 188728 172487 188730
rect 169894 188672 172426 188728
rect 172482 188672 172487 188728
rect 169894 188670 172487 188672
rect 169894 188360 169954 188670
rect 172421 188667 172487 188670
rect 303061 187642 303127 187645
rect 299828 187640 303127 187642
rect 299828 187584 303066 187640
rect 303122 187584 303127 187640
rect 299828 187582 303127 187584
rect 303061 187579 303127 187582
rect 172421 187370 172487 187373
rect 169894 187368 172487 187370
rect 169894 187312 172426 187368
rect 172482 187312 172487 187368
rect 169894 187310 172487 187312
rect 169894 187136 169954 187310
rect 172421 187307 172487 187310
rect 197353 187234 197419 187237
rect 197353 187232 200100 187234
rect 197353 187176 197358 187232
rect 197414 187176 200100 187232
rect 197353 187174 200100 187176
rect 197353 187171 197419 187174
rect 172421 186146 172487 186149
rect 169894 186144 172487 186146
rect 169894 186088 172426 186144
rect 172482 186088 172487 186144
rect 169894 186086 172487 186088
rect 169894 186048 169954 186086
rect 172421 186083 172487 186086
rect 198457 185194 198523 185197
rect 198457 185192 200100 185194
rect 198457 185136 198462 185192
rect 198518 185136 200100 185192
rect 198457 185134 200100 185136
rect 198457 185131 198523 185134
rect 169894 184786 169954 184824
rect 172421 184786 172487 184789
rect 169894 184784 172487 184786
rect 169894 184728 172426 184784
rect 172482 184728 172487 184784
rect 169894 184726 172487 184728
rect 172421 184723 172487 184726
rect 302785 184650 302851 184653
rect 299828 184648 302851 184650
rect 299828 184592 302790 184648
rect 302846 184592 302851 184648
rect 299828 184590 302851 184592
rect 302785 184587 302851 184590
rect 172329 184378 172395 184381
rect 169894 184376 172395 184378
rect 169894 184320 172334 184376
rect 172390 184320 172395 184376
rect 169894 184318 172395 184320
rect 169894 183736 169954 184318
rect 172329 184315 172395 184318
rect 172421 183018 172487 183021
rect 169894 183016 172487 183018
rect 169894 182960 172426 183016
rect 172482 182960 172487 183016
rect 169894 182958 172487 182960
rect 169894 182512 169954 182958
rect 172421 182955 172487 182958
rect 197353 183018 197419 183021
rect 197353 183016 200100 183018
rect 197353 182960 197358 183016
rect 197414 182960 200100 183016
rect 197353 182958 200100 182960
rect 197353 182955 197419 182958
rect 172421 181794 172487 181797
rect 169894 181792 172487 181794
rect 169894 181736 172426 181792
rect 172482 181736 172487 181792
rect 169894 181734 172487 181736
rect 169894 181424 169954 181734
rect 172421 181731 172487 181734
rect 302693 181522 302759 181525
rect 299828 181520 302759 181522
rect 299828 181464 302698 181520
rect 302754 181464 302759 181520
rect 299828 181462 302759 181464
rect 302693 181459 302759 181462
rect 198273 180978 198339 180981
rect 198273 180976 200100 180978
rect 198273 180920 198278 180976
rect 198334 180920 200100 180976
rect 198273 180918 200100 180920
rect 198273 180915 198339 180918
rect 172421 180570 172487 180573
rect 169894 180568 172487 180570
rect 169894 180512 172426 180568
rect 172482 180512 172487 180568
rect 169894 180510 172487 180512
rect 169894 180200 169954 180510
rect 172421 180507 172487 180510
rect 171133 179210 171199 179213
rect 169894 179208 171199 179210
rect 169894 179152 171138 179208
rect 171194 179152 171199 179208
rect 169894 179150 171199 179152
rect 169894 179112 169954 179150
rect 171133 179147 171199 179150
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 197353 178802 197419 178805
rect 197353 178800 200100 178802
rect 197353 178744 197358 178800
rect 197414 178744 200100 178800
rect 197353 178742 200100 178744
rect 197353 178739 197419 178742
rect 303337 178394 303403 178397
rect 299828 178392 303403 178394
rect 299828 178336 303342 178392
rect 303398 178336 303403 178392
rect 299828 178334 303403 178336
rect 303337 178331 303403 178334
rect 172421 177986 172487 177989
rect 169894 177984 172487 177986
rect 169894 177928 172426 177984
rect 172482 177928 172487 177984
rect 169894 177926 172487 177928
rect 169894 177888 169954 177926
rect 172421 177923 172487 177926
rect 172237 177442 172303 177445
rect 169894 177440 172303 177442
rect 169894 177384 172242 177440
rect 172298 177384 172303 177440
rect 169894 177382 172303 177384
rect 169894 176800 169954 177382
rect 172237 177379 172303 177382
rect 197353 176762 197419 176765
rect 197353 176760 200100 176762
rect 197353 176704 197358 176760
rect 197414 176704 200100 176760
rect 197353 176702 200100 176704
rect 197353 176699 197419 176702
rect 172237 176082 172303 176085
rect 169894 176080 172303 176082
rect -960 175796 480 176036
rect 169894 176024 172242 176080
rect 172298 176024 172303 176080
rect 169894 176022 172303 176024
rect 169894 175576 169954 176022
rect 172237 176019 172303 176022
rect 302233 175402 302299 175405
rect 299828 175400 302299 175402
rect 299828 175344 302238 175400
rect 302294 175344 302299 175400
rect 299828 175342 302299 175344
rect 302233 175339 302299 175342
rect 172421 174858 172487 174861
rect 169894 174856 172487 174858
rect 169894 174800 172426 174856
rect 172482 174800 172487 174856
rect 169894 174798 172487 174800
rect 169894 174488 169954 174798
rect 172421 174795 172487 174798
rect 197721 174586 197787 174589
rect 197721 174584 200100 174586
rect 197721 174528 197726 174584
rect 197782 174528 200100 174584
rect 197721 174526 200100 174528
rect 197721 174523 197787 174526
rect 172421 173634 172487 173637
rect 169894 173632 172487 173634
rect 169894 173576 172426 173632
rect 172482 173576 172487 173632
rect 169894 173574 172487 173576
rect 169894 173264 169954 173574
rect 172421 173571 172487 173574
rect 197353 172546 197419 172549
rect 197353 172544 200100 172546
rect 197353 172488 197358 172544
rect 197414 172488 200100 172544
rect 197353 172486 200100 172488
rect 197353 172483 197419 172486
rect 172421 172410 172487 172413
rect 169894 172408 172487 172410
rect 169894 172352 172426 172408
rect 172482 172352 172487 172408
rect 169894 172350 172487 172352
rect 169894 172176 169954 172350
rect 172421 172347 172487 172350
rect 303061 172274 303127 172277
rect 299828 172272 303127 172274
rect 299828 172216 303066 172272
rect 303122 172216 303127 172272
rect 299828 172214 303127 172216
rect 303061 172211 303127 172214
rect 172421 171050 172487 171053
rect 169894 171048 172487 171050
rect 169894 170992 172426 171048
rect 172482 170992 172487 171048
rect 169894 170990 172487 170992
rect 169894 170952 169954 170990
rect 172421 170987 172487 170990
rect 171777 170506 171843 170509
rect 169894 170504 171843 170506
rect 169894 170448 171782 170504
rect 171838 170448 171843 170504
rect 169894 170446 171843 170448
rect 169894 169864 169954 170446
rect 171777 170443 171843 170446
rect 197445 170370 197511 170373
rect 197445 170368 200100 170370
rect 197445 170312 197450 170368
rect 197506 170312 200100 170368
rect 197445 170310 200100 170312
rect 197445 170307 197511 170310
rect 444782 169628 444788 169692
rect 444852 169690 444858 169692
rect 445017 169690 445083 169693
rect 444852 169688 445083 169690
rect 444852 169632 445022 169688
rect 445078 169632 445083 169688
rect 444852 169630 445083 169632
rect 444852 169628 444858 169630
rect 445017 169627 445083 169630
rect 172237 169146 172303 169149
rect 302785 169146 302851 169149
rect 169894 169144 172303 169146
rect 169894 169088 172242 169144
rect 172298 169088 172303 169144
rect 169894 169086 172303 169088
rect 299828 169144 302851 169146
rect 299828 169088 302790 169144
rect 302846 169088 302851 169144
rect 299828 169086 302851 169088
rect 169894 168640 169954 169086
rect 172237 169083 172303 169086
rect 302785 169083 302851 169086
rect 372429 169010 372495 169013
rect 444782 169010 444788 169012
rect 372429 169008 444788 169010
rect 372429 168952 372434 169008
rect 372490 168952 444788 169008
rect 372429 168950 444788 168952
rect 372429 168947 372495 168950
rect 444782 168948 444788 168950
rect 444852 168948 444858 169012
rect 197353 168330 197419 168333
rect 197353 168328 200100 168330
rect 197353 168272 197358 168328
rect 197414 168272 200100 168328
rect 197353 168270 200100 168272
rect 197353 168267 197419 168270
rect 171869 168194 171935 168197
rect 169894 168192 171935 168194
rect 169894 168136 171874 168192
rect 171930 168136 171935 168192
rect 169894 168134 171935 168136
rect 169894 167552 169954 168134
rect 171869 168131 171935 168134
rect 172421 166698 172487 166701
rect 169894 166696 172487 166698
rect 169894 166640 172426 166696
rect 172482 166640 172487 166696
rect 169894 166638 172487 166640
rect 169894 166328 169954 166638
rect 172421 166635 172487 166638
rect 198457 166290 198523 166293
rect 198457 166288 200100 166290
rect 198457 166232 198462 166288
rect 198518 166232 200100 166288
rect 198457 166230 200100 166232
rect 198457 166227 198523 166230
rect 302785 166154 302851 166157
rect 299828 166152 302851 166154
rect 299828 166096 302790 166152
rect 302846 166096 302851 166152
rect 299828 166094 302851 166096
rect 302785 166091 302851 166094
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 169894 164522 169954 165240
rect 171961 164522 172027 164525
rect 169894 164520 172027 164522
rect 169894 164464 171966 164520
rect 172022 164464 172027 164520
rect 169894 164462 172027 164464
rect 171961 164459 172027 164462
rect 172053 164114 172119 164117
rect 169894 164112 172119 164114
rect 169894 164056 172058 164112
rect 172114 164056 172119 164112
rect 169894 164054 172119 164056
rect 169894 164016 169954 164054
rect 172053 164051 172119 164054
rect 197537 164114 197603 164117
rect 197537 164112 200100 164114
rect 197537 164056 197542 164112
rect 197598 164056 200100 164112
rect 197537 164054 200100 164056
rect 197537 164051 197603 164054
rect 172237 163570 172303 163573
rect 169894 163568 172303 163570
rect 169894 163512 172242 163568
rect 172298 163512 172303 163568
rect 169894 163510 172303 163512
rect -960 162890 480 162980
rect 169894 162928 169954 163510
rect 172237 163507 172303 163510
rect 302785 163026 302851 163029
rect 299828 163024 302851 163026
rect 299828 162968 302790 163024
rect 302846 162968 302851 163024
rect 299828 162966 302851 162968
rect 302785 162963 302851 162966
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 172145 162346 172211 162349
rect 169894 162344 172211 162346
rect 169894 162288 172150 162344
rect 172206 162288 172211 162344
rect 169894 162286 172211 162288
rect 169894 161704 169954 162286
rect 172145 162283 172211 162286
rect 198089 162074 198155 162077
rect 198089 162072 200100 162074
rect 198089 162016 198094 162072
rect 198150 162016 200100 162072
rect 198089 162014 200100 162016
rect 198089 162011 198155 162014
rect 172421 160986 172487 160989
rect 169894 160984 172487 160986
rect 169894 160928 172426 160984
rect 172482 160928 172487 160984
rect 169894 160926 172487 160928
rect 169894 160616 169954 160926
rect 172421 160923 172487 160926
rect 197537 159898 197603 159901
rect 302509 159898 302575 159901
rect 197537 159896 200100 159898
rect 197537 159840 197542 159896
rect 197598 159840 200100 159896
rect 197537 159838 200100 159840
rect 299828 159896 302575 159898
rect 299828 159840 302514 159896
rect 302570 159840 302575 159896
rect 299828 159838 302575 159840
rect 197537 159835 197603 159838
rect 302509 159835 302575 159838
rect 371918 158748 371924 158812
rect 371988 158810 371994 158812
rect 372153 158810 372219 158813
rect 442809 158810 442875 158813
rect 444598 158810 444604 158812
rect 371988 158808 444604 158810
rect 371988 158752 372158 158808
rect 372214 158752 442814 158808
rect 442870 158752 444604 158808
rect 371988 158750 444604 158752
rect 371988 158748 371994 158750
rect 372153 158747 372219 158750
rect 442809 158747 442875 158750
rect 444598 158748 444604 158750
rect 444668 158748 444674 158812
rect 197353 157858 197419 157861
rect 197353 157856 200100 157858
rect 197353 157800 197358 157856
rect 197414 157800 200100 157856
rect 197353 157798 200100 157800
rect 197353 157795 197419 157798
rect 302785 156906 302851 156909
rect 299828 156904 302851 156906
rect 299828 156848 302790 156904
rect 302846 156848 302851 156904
rect 299828 156846 302851 156848
rect 302785 156843 302851 156846
rect 444782 156436 444788 156500
rect 444852 156498 444858 156500
rect 445937 156498 446003 156501
rect 444852 156496 446003 156498
rect 444852 156440 445942 156496
rect 445998 156440 446003 156496
rect 444852 156438 446003 156440
rect 444852 156436 444858 156438
rect 445937 156435 446003 156438
rect 445937 156090 446003 156093
rect 513925 156090 513991 156093
rect 445937 156088 513991 156090
rect 445937 156032 445942 156088
rect 445998 156032 513930 156088
rect 513986 156032 513991 156088
rect 445937 156030 513991 156032
rect 445937 156027 446003 156030
rect 513925 156027 513991 156030
rect 197537 155682 197603 155685
rect 197537 155680 200100 155682
rect 197537 155624 197542 155680
rect 197598 155624 200100 155680
rect 197537 155622 200100 155624
rect 197537 155619 197603 155622
rect 441797 154050 441863 154053
rect 441797 154048 441906 154050
rect 441797 153992 441802 154048
rect 441858 153992 441906 154048
rect 441797 153987 441906 153992
rect 172329 153778 172395 153781
rect 302785 153778 302851 153781
rect 372102 153778 372108 153780
rect 169924 153776 172395 153778
rect 169924 153720 172334 153776
rect 172390 153720 172395 153776
rect 169924 153718 172395 153720
rect 299828 153776 302851 153778
rect 299828 153720 302790 153776
rect 302846 153720 302851 153776
rect 299828 153718 302851 153720
rect 369932 153718 372108 153778
rect 172329 153715 172395 153718
rect 302785 153715 302851 153718
rect 372102 153716 372108 153718
rect 372172 153716 372178 153780
rect 197353 153642 197419 153645
rect 197353 153640 200100 153642
rect 197353 153584 197358 153640
rect 197414 153584 200100 153640
rect 197353 153582 200100 153584
rect 197353 153579 197419 153582
rect 441846 153476 441906 153987
rect 483657 153914 483723 153917
rect 513557 153914 513623 153917
rect 483657 153912 513623 153914
rect 483657 153856 483662 153912
rect 483718 153856 513562 153912
rect 513618 153856 513623 153912
rect 483657 153854 513623 153856
rect 483657 153851 483723 153854
rect 513557 153851 513623 153854
rect 516869 153778 516935 153781
rect 513820 153776 516935 153778
rect 513820 153720 516874 153776
rect 516930 153720 516935 153776
rect 513820 153718 516935 153720
rect 516869 153715 516935 153718
rect 172237 153234 172303 153237
rect 372286 153234 372292 153236
rect 169924 153232 172303 153234
rect 169924 153176 172242 153232
rect 172298 153176 172303 153232
rect 169924 153174 172303 153176
rect 369932 153174 372292 153234
rect 172237 153171 172303 153174
rect 372286 153172 372292 153174
rect 372356 153172 372362 153236
rect 517605 153234 517671 153237
rect 513820 153232 517671 153234
rect 513820 153176 517610 153232
rect 517666 153176 517671 153232
rect 513820 153174 517671 153176
rect 517605 153171 517671 153174
rect 371233 152964 371299 152965
rect 371182 152900 371188 152964
rect 371252 152962 371299 152964
rect 513373 152962 513439 152965
rect 514150 152962 514156 152964
rect 371252 152960 371344 152962
rect 371294 152904 371344 152960
rect 371252 152902 371344 152904
rect 513373 152960 514156 152962
rect 513373 152904 513378 152960
rect 513434 152904 514156 152960
rect 513373 152902 514156 152904
rect 371252 152900 371299 152902
rect 371233 152899 371299 152900
rect 513373 152899 513439 152902
rect 514150 152900 514156 152902
rect 514220 152900 514226 152964
rect 172421 152690 172487 152693
rect 371550 152690 371556 152692
rect 169924 152688 172487 152690
rect 169924 152632 172426 152688
rect 172482 152632 172487 152688
rect 169924 152630 172487 152632
rect 369932 152630 371556 152690
rect 172421 152627 172487 152630
rect 371550 152628 371556 152630
rect 371620 152628 371626 152692
rect 516133 152690 516199 152693
rect 513820 152688 516199 152690
rect 513820 152632 516138 152688
rect 516194 152632 516199 152688
rect 513820 152630 516199 152632
rect 516133 152627 516199 152630
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 445661 152418 445727 152421
rect 441876 152416 445727 152418
rect 441876 152388 445666 152416
rect 441846 152360 445666 152388
rect 445722 152360 445727 152416
rect 441846 152358 445727 152360
rect 172329 152146 172395 152149
rect 371734 152146 371740 152148
rect 169924 152144 172395 152146
rect 169924 152088 172334 152144
rect 172390 152088 172395 152144
rect 169924 152086 172395 152088
rect 369932 152086 371740 152146
rect 172329 152083 172395 152086
rect 371734 152084 371740 152086
rect 371804 152084 371810 152148
rect 441846 152013 441906 152358
rect 445661 152355 445727 152358
rect 513833 152418 513899 152421
rect 513966 152418 513972 152420
rect 513833 152416 513972 152418
rect 513833 152360 513838 152416
rect 513894 152360 513972 152416
rect 513833 152358 513972 152360
rect 513833 152355 513899 152358
rect 513966 152356 513972 152358
rect 514036 152356 514042 152420
rect 516225 152146 516291 152149
rect 513820 152144 516291 152146
rect 513820 152088 516230 152144
rect 516286 152088 516291 152144
rect 513820 152086 516291 152088
rect 516225 152083 516291 152086
rect 441797 152008 441906 152013
rect 514385 152012 514451 152013
rect 441797 151952 441802 152008
rect 441858 151952 441906 152008
rect 441797 151950 441906 151952
rect 441797 151947 441863 151950
rect 514334 151948 514340 152012
rect 514404 152010 514451 152012
rect 514404 152008 514496 152010
rect 514446 151952 514496 152008
rect 514404 151950 514496 151952
rect 514404 151948 514451 151950
rect 514385 151947 514451 151948
rect 514150 151812 514156 151876
rect 514220 151874 514226 151876
rect 514385 151874 514451 151877
rect 514220 151872 514451 151874
rect 514220 151816 514390 151872
rect 514446 151816 514451 151872
rect 514220 151814 514451 151816
rect 514220 151812 514226 151814
rect 514385 151811 514451 151814
rect 369301 151738 369367 151741
rect 513557 151738 513623 151741
rect 369301 151736 369410 151738
rect 369301 151680 369306 151736
rect 369362 151680 369410 151736
rect 369301 151675 369410 151680
rect 513557 151736 513666 151738
rect 513557 151680 513562 151736
rect 513618 151680 513666 151736
rect 513557 151675 513666 151680
rect 171685 151602 171751 151605
rect 169924 151600 171751 151602
rect 169924 151544 171690 151600
rect 171746 151544 171751 151600
rect 369350 151572 369410 151675
rect 513606 151572 513666 151675
rect 169924 151542 171751 151544
rect 171685 151539 171751 151542
rect 197537 151466 197603 151469
rect 514201 151466 514267 151469
rect 514334 151466 514340 151468
rect 197537 151464 200100 151466
rect 197537 151408 197542 151464
rect 197598 151408 200100 151464
rect 197537 151406 200100 151408
rect 514201 151464 514340 151466
rect 514201 151408 514206 151464
rect 514262 151408 514340 151464
rect 514201 151406 514340 151408
rect 197537 151403 197603 151406
rect 514201 151403 514267 151406
rect 514334 151404 514340 151406
rect 514404 151404 514410 151468
rect 369485 151330 369551 151333
rect 513649 151330 513715 151333
rect 369485 151328 369594 151330
rect 369485 151272 369490 151328
rect 369546 151272 369594 151328
rect 369485 151267 369594 151272
rect 171501 151058 171567 151061
rect 169924 151056 171567 151058
rect 169924 151000 171506 151056
rect 171562 151000 171567 151056
rect 369534 151028 369594 151267
rect 513606 151328 513715 151330
rect 513606 151272 513654 151328
rect 513710 151272 513715 151328
rect 513606 151267 513715 151272
rect 513966 151268 513972 151332
rect 514036 151330 514042 151332
rect 514109 151330 514175 151333
rect 514036 151328 514175 151330
rect 514036 151272 514114 151328
rect 514170 151272 514175 151328
rect 514036 151270 514175 151272
rect 514036 151268 514042 151270
rect 514109 151267 514175 151270
rect 445937 151194 446003 151197
rect 441876 151192 446003 151194
rect 441876 151136 445942 151192
rect 445998 151136 446003 151192
rect 441876 151134 446003 151136
rect 445937 151131 446003 151134
rect 513606 151028 513666 151267
rect 169924 150998 171567 151000
rect 171501 150995 171567 150998
rect 302785 150786 302851 150789
rect 369577 150786 369643 150789
rect 514293 150786 514359 150789
rect 299828 150784 302851 150786
rect 299828 150728 302790 150784
rect 302846 150728 302851 150784
rect 299828 150726 302851 150728
rect 302785 150723 302851 150726
rect 369534 150784 369643 150786
rect 369534 150728 369582 150784
rect 369638 150728 369643 150784
rect 369534 150723 369643 150728
rect 513790 150784 514359 150786
rect 513790 150728 514298 150784
rect 514354 150728 514359 150784
rect 513790 150726 514359 150728
rect 171593 150514 171659 150517
rect 169924 150512 171659 150514
rect 169924 150456 171598 150512
rect 171654 150456 171659 150512
rect 369534 150484 369594 150723
rect 513790 150484 513850 150726
rect 514293 150723 514359 150726
rect 169924 150454 171659 150456
rect 171593 150451 171659 150454
rect 442717 150378 442783 150381
rect 441846 150376 442783 150378
rect 441846 150320 442722 150376
rect 442778 150320 442783 150376
rect 441846 150318 442783 150320
rect 441846 150076 441906 150318
rect 442717 150315 442783 150318
rect 513741 150242 513807 150245
rect 513741 150240 513850 150242
rect 513741 150184 513746 150240
rect 513802 150184 513850 150240
rect 513741 150179 513850 150184
rect 171685 149970 171751 149973
rect 370405 149970 370471 149973
rect 169924 149968 171751 149970
rect -960 149834 480 149924
rect 169924 149912 171690 149968
rect 171746 149912 171751 149968
rect 169924 149910 171751 149912
rect 369932 149968 370471 149970
rect 369932 149912 370410 149968
rect 370466 149912 370471 149968
rect 513790 149940 513850 150179
rect 369932 149910 370471 149912
rect 171685 149907 171751 149910
rect 370405 149907 370471 149910
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 513373 149698 513439 149701
rect 513373 149696 513482 149698
rect 513373 149640 513378 149696
rect 513434 149640 513482 149696
rect 513373 149635 513482 149640
rect 171685 149426 171751 149429
rect 169924 149424 171751 149426
rect 169924 149368 171690 149424
rect 171746 149368 171751 149424
rect 169924 149366 171751 149368
rect 171685 149363 171751 149366
rect 197353 149426 197419 149429
rect 371233 149426 371299 149429
rect 197353 149424 200100 149426
rect 197353 149368 197358 149424
rect 197414 149368 200100 149424
rect 197353 149366 200100 149368
rect 369932 149424 371299 149426
rect 369932 149368 371238 149424
rect 371294 149368 371299 149424
rect 513422 149396 513482 149635
rect 369932 149366 371299 149368
rect 197353 149363 197419 149366
rect 371233 149363 371299 149366
rect 513281 149018 513347 149021
rect 513281 149016 513482 149018
rect 513281 148960 513286 149016
rect 513342 148960 513482 149016
rect 513281 148958 513482 148960
rect 513281 148955 513347 148958
rect 172237 148882 172303 148885
rect 370313 148882 370379 148885
rect 445293 148882 445359 148885
rect 169924 148880 172303 148882
rect 169924 148824 172242 148880
rect 172298 148824 172303 148880
rect 169924 148822 172303 148824
rect 369932 148880 370379 148882
rect 369932 148824 370318 148880
rect 370374 148824 370379 148880
rect 369932 148822 370379 148824
rect 441876 148880 445359 148882
rect 441876 148824 445298 148880
rect 445354 148824 445359 148880
rect 513422 148852 513482 148958
rect 441876 148822 445359 148824
rect 172237 148819 172303 148822
rect 370313 148819 370379 148822
rect 445293 148819 445359 148822
rect 513465 148610 513531 148613
rect 513422 148608 513531 148610
rect 513422 148552 513470 148608
rect 513526 148552 513531 148608
rect 513422 148547 513531 148552
rect 171685 148338 171751 148341
rect 371182 148338 371188 148340
rect 169924 148336 171751 148338
rect 169924 148280 171690 148336
rect 171746 148280 171751 148336
rect 169924 148278 171751 148280
rect 369932 148278 371188 148338
rect 171685 148275 171751 148278
rect 371182 148276 371188 148278
rect 371252 148276 371258 148340
rect 513422 148308 513482 148547
rect 171501 147794 171567 147797
rect 371325 147794 371391 147797
rect 444373 147794 444439 147797
rect 516317 147794 516383 147797
rect 169924 147792 171567 147794
rect 169924 147736 171506 147792
rect 171562 147736 171567 147792
rect 169924 147734 171567 147736
rect 369932 147792 371391 147794
rect 369932 147736 371330 147792
rect 371386 147736 371391 147792
rect 369932 147734 371391 147736
rect 441876 147792 444439 147794
rect 441876 147736 444378 147792
rect 444434 147736 444439 147792
rect 441876 147734 444439 147736
rect 513820 147792 516383 147794
rect 513820 147736 516322 147792
rect 516378 147736 516383 147792
rect 513820 147734 516383 147736
rect 171501 147731 171567 147734
rect 371325 147731 371391 147734
rect 444373 147731 444439 147734
rect 516317 147731 516383 147734
rect 302693 147658 302759 147661
rect 299828 147656 302759 147658
rect 299828 147600 302698 147656
rect 302754 147600 302759 147656
rect 299828 147598 302759 147600
rect 302693 147595 302759 147598
rect 172421 147250 172487 147253
rect 169924 147248 172487 147250
rect 169924 147192 172426 147248
rect 172482 147192 172487 147248
rect 169924 147190 172487 147192
rect 172421 147187 172487 147190
rect 197629 147250 197695 147253
rect 371325 147250 371391 147253
rect 516225 147250 516291 147253
rect 197629 147248 200100 147250
rect 197629 147192 197634 147248
rect 197690 147192 200100 147248
rect 197629 147190 200100 147192
rect 369932 147248 371391 147250
rect 369932 147192 371330 147248
rect 371386 147192 371391 147248
rect 369932 147190 371391 147192
rect 513820 147248 516291 147250
rect 513820 147192 516230 147248
rect 516286 147192 516291 147248
rect 513820 147190 516291 147192
rect 197629 147187 197695 147190
rect 371325 147187 371391 147190
rect 516225 147187 516291 147190
rect 171501 146706 171567 146709
rect 371969 146706 372035 146709
rect 516685 146706 516751 146709
rect 169924 146704 171567 146706
rect 169924 146648 171506 146704
rect 171562 146648 171567 146704
rect 169924 146646 171567 146648
rect 369932 146704 372035 146706
rect 369932 146648 371974 146704
rect 372030 146648 372035 146704
rect 369932 146646 372035 146648
rect 513820 146704 516751 146706
rect 513820 146648 516690 146704
rect 516746 146648 516751 146704
rect 513820 146646 516751 146648
rect 171501 146643 171567 146646
rect 371969 146643 372035 146646
rect 516685 146643 516751 146646
rect 443085 146570 443151 146573
rect 441876 146568 443151 146570
rect 441876 146512 443090 146568
rect 443146 146512 443151 146568
rect 441876 146510 443151 146512
rect 443085 146507 443151 146510
rect 172329 146162 172395 146165
rect 371969 146162 372035 146165
rect 514293 146162 514359 146165
rect 169924 146160 172395 146162
rect 169924 146104 172334 146160
rect 172390 146104 172395 146160
rect 169924 146102 172395 146104
rect 369932 146160 372035 146162
rect 369932 146104 371974 146160
rect 372030 146104 372035 146160
rect 369932 146102 372035 146104
rect 513820 146160 514359 146162
rect 513820 146104 514298 146160
rect 514354 146104 514359 146160
rect 513820 146102 514359 146104
rect 172329 146099 172395 146102
rect 371969 146099 372035 146102
rect 514293 146099 514359 146102
rect 442257 146026 442323 146029
rect 441846 146024 442323 146026
rect 441846 145968 442262 146024
rect 442318 145968 442323 146024
rect 441846 145966 442323 145968
rect 172421 145618 172487 145621
rect 371325 145618 371391 145621
rect 169924 145616 172487 145618
rect 169924 145560 172426 145616
rect 172482 145560 172487 145616
rect 169924 145558 172487 145560
rect 369932 145616 371391 145618
rect 369932 145560 371330 145616
rect 371386 145560 371391 145616
rect 369932 145558 371391 145560
rect 172421 145555 172487 145558
rect 371325 145555 371391 145558
rect 441846 145452 441906 145966
rect 442257 145963 442323 145966
rect 516133 145618 516199 145621
rect 513820 145616 516199 145618
rect 513820 145560 516138 145616
rect 516194 145560 516199 145616
rect 513820 145558 516199 145560
rect 516133 145555 516199 145558
rect 197353 145210 197419 145213
rect 197353 145208 200100 145210
rect 197353 145152 197358 145208
rect 197414 145152 200100 145208
rect 197353 145150 200100 145152
rect 197353 145147 197419 145150
rect 171501 145074 171567 145077
rect 371325 145074 371391 145077
rect 516409 145074 516475 145077
rect 169924 145072 171567 145074
rect 169924 145016 171506 145072
rect 171562 145016 171567 145072
rect 169924 145014 171567 145016
rect 369932 145072 371391 145074
rect 369932 145016 371330 145072
rect 371386 145016 371391 145072
rect 369932 145014 371391 145016
rect 513820 145072 516475 145074
rect 513820 145016 516414 145072
rect 516470 145016 516475 145072
rect 513820 145014 516475 145016
rect 171501 145011 171567 145014
rect 371325 145011 371391 145014
rect 516409 145011 516475 145014
rect 172421 144530 172487 144533
rect 302785 144530 302851 144533
rect 371325 144530 371391 144533
rect 516593 144530 516659 144533
rect 169924 144528 172487 144530
rect 169924 144472 172426 144528
rect 172482 144472 172487 144528
rect 169924 144470 172487 144472
rect 299828 144528 302851 144530
rect 299828 144472 302790 144528
rect 302846 144472 302851 144528
rect 299828 144470 302851 144472
rect 369932 144528 371391 144530
rect 369932 144472 371330 144528
rect 371386 144472 371391 144528
rect 369932 144470 371391 144472
rect 513820 144528 516659 144530
rect 513820 144472 516598 144528
rect 516654 144472 516659 144528
rect 513820 144470 516659 144472
rect 172421 144467 172487 144470
rect 302785 144467 302851 144470
rect 371325 144467 371391 144470
rect 516593 144467 516659 144470
rect 444833 144258 444899 144261
rect 441876 144256 444899 144258
rect 441876 144200 444838 144256
rect 444894 144200 444899 144256
rect 441876 144198 444899 144200
rect 444833 144195 444899 144198
rect 171777 144122 171843 144125
rect 371325 144122 371391 144125
rect 516777 144122 516843 144125
rect 169924 144120 171843 144122
rect 169924 144064 171782 144120
rect 171838 144064 171843 144120
rect 169924 144062 171843 144064
rect 369932 144120 371391 144122
rect 369932 144064 371330 144120
rect 371386 144064 371391 144120
rect 369932 144062 371391 144064
rect 513820 144120 516843 144122
rect 513820 144064 516782 144120
rect 516838 144064 516843 144120
rect 513820 144062 516843 144064
rect 171777 144059 171843 144062
rect 371325 144059 371391 144062
rect 516777 144059 516843 144062
rect 369393 143850 369459 143853
rect 369350 143848 369459 143850
rect 369350 143792 369398 143848
rect 369454 143792 369459 143848
rect 369350 143787 369459 143792
rect 171961 143578 172027 143581
rect 169924 143576 172027 143578
rect 169924 143520 171966 143576
rect 172022 143520 172027 143576
rect 369350 143548 369410 143787
rect 516501 143578 516567 143581
rect 513820 143576 516567 143578
rect 169924 143518 172027 143520
rect 513820 143520 516506 143576
rect 516562 143520 516567 143576
rect 513820 143518 516567 143520
rect 171961 143515 172027 143518
rect 516501 143515 516567 143518
rect 445109 143170 445175 143173
rect 441876 143168 445175 143170
rect 441876 143112 445114 143168
rect 445170 143112 445175 143168
rect 441876 143110 445175 143112
rect 445109 143107 445175 143110
rect 172237 143034 172303 143037
rect 169924 143032 172303 143034
rect 169924 142976 172242 143032
rect 172298 142976 172303 143032
rect 169924 142974 172303 142976
rect 172237 142971 172303 142974
rect 197353 143034 197419 143037
rect 371969 143034 372035 143037
rect 515581 143034 515647 143037
rect 197353 143032 200100 143034
rect 197353 142976 197358 143032
rect 197414 142976 200100 143032
rect 197353 142974 200100 142976
rect 369932 143032 372035 143034
rect 369932 142976 371974 143032
rect 372030 142976 372035 143032
rect 369932 142974 372035 142976
rect 513820 143032 515647 143034
rect 513820 142976 515586 143032
rect 515642 142976 515647 143032
rect 513820 142974 515647 142976
rect 197353 142971 197419 142974
rect 371969 142971 372035 142974
rect 515581 142971 515647 142974
rect 513281 142762 513347 142765
rect 513281 142760 513482 142762
rect 513281 142704 513286 142760
rect 513342 142704 513482 142760
rect 513281 142702 513482 142704
rect 513281 142699 513347 142702
rect 171593 142490 171659 142493
rect 371325 142490 371391 142493
rect 169924 142488 171659 142490
rect 169924 142432 171598 142488
rect 171654 142432 171659 142488
rect 169924 142430 171659 142432
rect 369932 142488 371391 142490
rect 369932 142432 371330 142488
rect 371386 142432 371391 142488
rect 513422 142460 513482 142702
rect 369932 142430 371391 142432
rect 171593 142427 171659 142430
rect 371325 142427 371391 142430
rect 171409 141946 171475 141949
rect 370221 141946 370287 141949
rect 445201 141946 445267 141949
rect 515213 141946 515279 141949
rect 169924 141944 171475 141946
rect 169924 141888 171414 141944
rect 171470 141888 171475 141944
rect 169924 141886 171475 141888
rect 369932 141944 370287 141946
rect 369932 141888 370226 141944
rect 370282 141888 370287 141944
rect 369932 141886 370287 141888
rect 441876 141944 445267 141946
rect 441876 141888 445206 141944
rect 445262 141888 445267 141944
rect 441876 141886 445267 141888
rect 513820 141944 515279 141946
rect 513820 141888 515218 141944
rect 515274 141888 515279 141944
rect 513820 141886 515279 141888
rect 171409 141883 171475 141886
rect 370221 141883 370287 141886
rect 445201 141883 445267 141886
rect 515213 141883 515279 141886
rect 302325 141538 302391 141541
rect 299828 141536 302391 141538
rect 299828 141480 302330 141536
rect 302386 141480 302391 141536
rect 299828 141478 302391 141480
rect 302325 141475 302391 141478
rect 171501 141402 171567 141405
rect 371969 141402 372035 141405
rect 514293 141402 514359 141405
rect 169924 141400 171567 141402
rect 169924 141344 171506 141400
rect 171562 141344 171567 141400
rect 169924 141342 171567 141344
rect 369932 141400 372035 141402
rect 369932 141344 371974 141400
rect 372030 141344 372035 141400
rect 369932 141342 372035 141344
rect 513820 141400 514359 141402
rect 513820 141344 514298 141400
rect 514354 141344 514359 141400
rect 513820 141342 514359 141344
rect 171501 141339 171567 141342
rect 371969 141339 372035 141342
rect 514293 141339 514359 141342
rect 197353 140994 197419 140997
rect 197353 140992 200100 140994
rect 197353 140936 197358 140992
rect 197414 140936 200100 140992
rect 197353 140934 200100 140936
rect 197353 140931 197419 140934
rect 172421 140858 172487 140861
rect 370589 140858 370655 140861
rect 444649 140858 444715 140861
rect 515121 140858 515187 140861
rect 169924 140856 172487 140858
rect 169924 140800 172426 140856
rect 172482 140800 172487 140856
rect 169924 140798 172487 140800
rect 369932 140856 370655 140858
rect 369932 140800 370594 140856
rect 370650 140800 370655 140856
rect 369932 140798 370655 140800
rect 441876 140856 444715 140858
rect 441876 140800 444654 140856
rect 444710 140800 444715 140856
rect 441876 140798 444715 140800
rect 513820 140856 515187 140858
rect 513820 140800 515126 140856
rect 515182 140800 515187 140856
rect 513820 140798 515187 140800
rect 172421 140795 172487 140798
rect 370589 140795 370655 140798
rect 444649 140795 444715 140798
rect 515121 140795 515187 140798
rect 171501 140314 171567 140317
rect 370497 140314 370563 140317
rect 515029 140314 515095 140317
rect 169924 140312 171567 140314
rect 169924 140256 171506 140312
rect 171562 140256 171567 140312
rect 169924 140254 171567 140256
rect 369932 140312 370563 140314
rect 369932 140256 370502 140312
rect 370558 140256 370563 140312
rect 369932 140254 370563 140256
rect 513820 140312 515095 140314
rect 513820 140256 515034 140312
rect 515090 140256 515095 140312
rect 513820 140254 515095 140256
rect 171501 140251 171567 140254
rect 370497 140251 370563 140254
rect 515029 140251 515095 140254
rect 171685 139770 171751 139773
rect 370129 139770 370195 139773
rect 515305 139770 515371 139773
rect 169924 139768 171751 139770
rect 169924 139712 171690 139768
rect 171746 139712 171751 139768
rect 169924 139710 171751 139712
rect 369932 139768 370195 139770
rect 369932 139712 370134 139768
rect 370190 139712 370195 139768
rect 369932 139710 370195 139712
rect 513820 139768 515371 139770
rect 513820 139712 515310 139768
rect 515366 139712 515371 139768
rect 513820 139710 515371 139712
rect 171685 139707 171751 139710
rect 370129 139707 370195 139710
rect 515305 139707 515371 139710
rect 445569 139634 445635 139637
rect 441876 139632 445635 139634
rect 441876 139576 445574 139632
rect 445630 139576 445635 139632
rect 441876 139574 445635 139576
rect 445569 139571 445635 139574
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 172421 139226 172487 139229
rect 372153 139226 372219 139229
rect 515489 139226 515555 139229
rect 169924 139224 172487 139226
rect 169924 139168 172426 139224
rect 172482 139168 172487 139224
rect 169924 139166 172487 139168
rect 369932 139224 372219 139226
rect 369932 139168 372158 139224
rect 372214 139168 372219 139224
rect 369932 139166 372219 139168
rect 513820 139224 515555 139226
rect 513820 139168 515494 139224
rect 515550 139168 515555 139224
rect 583520 139212 584960 139302
rect 513820 139166 515555 139168
rect 172421 139163 172487 139166
rect 372153 139163 372219 139166
rect 515489 139163 515555 139166
rect 197353 138818 197419 138821
rect 197353 138816 200100 138818
rect 197353 138760 197358 138816
rect 197414 138760 200100 138816
rect 197353 138758 200100 138760
rect 197353 138755 197419 138758
rect 171869 138682 171935 138685
rect 371693 138682 371759 138685
rect 516501 138682 516567 138685
rect 169924 138680 171935 138682
rect 169924 138624 171874 138680
rect 171930 138624 171935 138680
rect 169924 138622 171935 138624
rect 369932 138680 371759 138682
rect 369932 138624 371698 138680
rect 371754 138624 371759 138680
rect 369932 138622 371759 138624
rect 513820 138680 516567 138682
rect 513820 138624 516506 138680
rect 516562 138624 516567 138680
rect 513820 138622 516567 138624
rect 171869 138619 171935 138622
rect 371693 138619 371759 138622
rect 516501 138619 516567 138622
rect 445845 138546 445911 138549
rect 441876 138544 445911 138546
rect 441876 138488 445850 138544
rect 445906 138488 445911 138544
rect 441876 138486 445911 138488
rect 445845 138483 445911 138486
rect 302877 138410 302943 138413
rect 299828 138408 302943 138410
rect 299828 138352 302882 138408
rect 302938 138352 302943 138408
rect 299828 138350 302943 138352
rect 302877 138347 302943 138350
rect 171685 138138 171751 138141
rect 371325 138138 371391 138141
rect 516225 138138 516291 138141
rect 169924 138136 171751 138138
rect 169924 138080 171690 138136
rect 171746 138080 171751 138136
rect 169924 138078 171751 138080
rect 369932 138136 371391 138138
rect 369932 138080 371330 138136
rect 371386 138080 371391 138136
rect 369932 138078 371391 138080
rect 513820 138136 516291 138138
rect 513820 138080 516230 138136
rect 516286 138080 516291 138136
rect 513820 138078 516291 138080
rect 171685 138075 171751 138078
rect 371325 138075 371391 138078
rect 516225 138075 516291 138078
rect 172421 137594 172487 137597
rect 371325 137594 371391 137597
rect 516133 137594 516199 137597
rect 169924 137592 172487 137594
rect 169924 137536 172426 137592
rect 172482 137536 172487 137592
rect 169924 137534 172487 137536
rect 369932 137592 371391 137594
rect 369932 137536 371330 137592
rect 371386 137536 371391 137592
rect 369932 137534 371391 137536
rect 513820 137592 516199 137594
rect 513820 137536 516138 137592
rect 516194 137536 516199 137592
rect 513820 137534 516199 137536
rect 172421 137531 172487 137534
rect 371325 137531 371391 137534
rect 516133 137531 516199 137534
rect 442993 137322 443059 137325
rect 445293 137322 445359 137325
rect 513925 137322 513991 137325
rect 441876 137320 445359 137322
rect 441876 137264 442998 137320
rect 443054 137264 445298 137320
rect 445354 137264 445359 137320
rect 441876 137262 445359 137264
rect 442993 137259 443059 137262
rect 445293 137259 445359 137262
rect 513790 137320 513991 137322
rect 513790 137264 513930 137320
rect 513986 137264 513991 137320
rect 513790 137262 513991 137264
rect 172237 137050 172303 137053
rect 372797 137050 372863 137053
rect 169924 137048 172303 137050
rect 169924 136992 172242 137048
rect 172298 136992 172303 137048
rect 169924 136990 172303 136992
rect 369932 137048 372863 137050
rect 369932 136992 372802 137048
rect 372858 136992 372863 137048
rect 513790 137020 513850 137262
rect 513925 137259 513991 137262
rect 369932 136990 372863 136992
rect 172237 136987 172303 136990
rect 372797 136987 372863 136990
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 197353 136778 197419 136781
rect 197353 136776 200100 136778
rect 197353 136720 197358 136776
rect 197414 136720 200100 136776
rect 197353 136718 200100 136720
rect 197353 136715 197419 136718
rect 369301 136642 369367 136645
rect 513833 136642 513899 136645
rect 369301 136640 369410 136642
rect 369301 136584 369306 136640
rect 369362 136584 369410 136640
rect 369301 136579 369410 136584
rect 172329 136506 172395 136509
rect 169924 136504 172395 136506
rect 169924 136448 172334 136504
rect 172390 136448 172395 136504
rect 369350 136476 369410 136579
rect 513790 136640 513899 136642
rect 513790 136584 513838 136640
rect 513894 136584 513899 136640
rect 513790 136579 513899 136584
rect 513790 136476 513850 136579
rect 169924 136446 172395 136448
rect 172329 136443 172395 136446
rect 441662 135965 441722 136204
rect 172421 135962 172487 135965
rect 371969 135962 372035 135965
rect 169924 135960 172487 135962
rect 169924 135904 172426 135960
rect 172482 135904 172487 135960
rect 169924 135902 172487 135904
rect 369932 135960 372035 135962
rect 369932 135904 371974 135960
rect 372030 135904 372035 135960
rect 369932 135902 372035 135904
rect 172421 135899 172487 135902
rect 371969 135899 372035 135902
rect 441613 135960 441722 135965
rect 514937 135962 515003 135965
rect 441613 135904 441618 135960
rect 441674 135904 441722 135960
rect 441613 135902 441722 135904
rect 513820 135960 515003 135962
rect 513820 135904 514942 135960
rect 514998 135904 515003 135960
rect 513820 135902 515003 135904
rect 441613 135899 441679 135902
rect 514937 135899 515003 135902
rect 172237 135418 172303 135421
rect 372337 135418 372403 135421
rect 514201 135418 514267 135421
rect 169924 135416 172303 135418
rect 169924 135360 172242 135416
rect 172298 135360 172303 135416
rect 169924 135358 172303 135360
rect 369932 135416 372403 135418
rect 369932 135360 372342 135416
rect 372398 135360 372403 135416
rect 369932 135358 372403 135360
rect 513820 135416 514267 135418
rect 513820 135360 514206 135416
rect 514262 135360 514267 135416
rect 513820 135358 514267 135360
rect 172237 135355 172303 135358
rect 372337 135355 372403 135358
rect 514201 135355 514267 135358
rect 302969 135282 303035 135285
rect 299828 135280 303035 135282
rect 299828 135224 302974 135280
rect 303030 135224 303035 135280
rect 299828 135222 303035 135224
rect 302969 135219 303035 135222
rect 369301 135010 369367 135013
rect 443085 135010 443151 135013
rect 444414 135010 444420 135012
rect 369301 135008 369410 135010
rect 369301 134952 369306 135008
rect 369362 134952 369410 135008
rect 369301 134947 369410 134952
rect 441876 135008 444420 135010
rect 441876 134952 443090 135008
rect 443146 134952 444420 135008
rect 441876 134950 444420 134952
rect 443085 134947 443151 134950
rect 444414 134948 444420 134950
rect 444484 134948 444490 135012
rect 172237 134874 172303 134877
rect 169924 134872 172303 134874
rect 169924 134816 172242 134872
rect 172298 134816 172303 134872
rect 369350 134844 369410 134947
rect 514845 134874 514911 134877
rect 513820 134872 514911 134874
rect 169924 134814 172303 134816
rect 513820 134816 514850 134872
rect 514906 134816 514911 134872
rect 513820 134814 514911 134816
rect 172237 134811 172303 134814
rect 514845 134811 514911 134814
rect 197721 134602 197787 134605
rect 197721 134600 200100 134602
rect 197721 134544 197726 134600
rect 197782 134544 200100 134600
rect 197721 134542 200100 134544
rect 197721 134539 197787 134542
rect 171869 134330 171935 134333
rect 371693 134330 371759 134333
rect 514753 134330 514819 134333
rect 169924 134328 171935 134330
rect 169924 134272 171874 134328
rect 171930 134272 171935 134328
rect 169924 134270 171935 134272
rect 369932 134328 371759 134330
rect 369932 134272 371698 134328
rect 371754 134272 371759 134328
rect 369932 134270 371759 134272
rect 513820 134328 514819 134330
rect 513820 134272 514758 134328
rect 514814 134272 514819 134328
rect 513820 134270 514819 134272
rect 171869 134267 171935 134270
rect 371693 134267 371759 134270
rect 514753 134267 514819 134270
rect 513373 134058 513439 134061
rect 513373 134056 513482 134058
rect 513373 134000 513378 134056
rect 513434 134000 513482 134056
rect 513373 133995 513482 134000
rect 171685 133922 171751 133925
rect 372521 133922 372587 133925
rect 445661 133922 445727 133925
rect 169924 133920 171751 133922
rect 169924 133864 171690 133920
rect 171746 133864 171751 133920
rect 169924 133862 171751 133864
rect 369932 133920 372587 133922
rect 369932 133864 372526 133920
rect 372582 133864 372587 133920
rect 369932 133862 372587 133864
rect 441876 133920 445727 133922
rect 441876 133864 445666 133920
rect 445722 133864 445727 133920
rect 513422 133892 513482 133995
rect 441876 133862 445727 133864
rect 171685 133859 171751 133862
rect 372521 133859 372587 133862
rect 445661 133859 445727 133862
rect 370037 133650 370103 133653
rect 513649 133650 513715 133653
rect 369902 133648 370103 133650
rect 369902 133592 370042 133648
rect 370098 133592 370103 133648
rect 369902 133590 370103 133592
rect 172513 133378 172579 133381
rect 169924 133376 172579 133378
rect 169924 133320 172518 133376
rect 172574 133320 172579 133376
rect 369902 133348 369962 133590
rect 370037 133587 370103 133590
rect 513606 133648 513715 133650
rect 513606 133592 513654 133648
rect 513710 133592 513715 133648
rect 513606 133587 513715 133592
rect 513606 133348 513666 133587
rect 169924 133318 172579 133320
rect 172513 133315 172579 133318
rect 513741 133106 513807 133109
rect 513741 133104 513850 133106
rect 513741 133048 513746 133104
rect 513802 133048 513850 133104
rect 513741 133043 513850 133048
rect 172421 132834 172487 132837
rect 371509 132834 371575 132837
rect 169924 132832 172487 132834
rect 169924 132776 172426 132832
rect 172482 132776 172487 132832
rect 169924 132774 172487 132776
rect 369932 132832 371575 132834
rect 369932 132776 371514 132832
rect 371570 132776 371575 132832
rect 513790 132804 513850 133043
rect 369932 132774 371575 132776
rect 172421 132771 172487 132774
rect 371509 132771 371575 132774
rect 445109 132698 445175 132701
rect 441876 132696 445175 132698
rect 441876 132640 445114 132696
rect 445170 132640 445175 132696
rect 441876 132638 445175 132640
rect 445109 132635 445175 132638
rect 197353 132562 197419 132565
rect 197353 132560 200100 132562
rect 197353 132504 197358 132560
rect 197414 132504 200100 132560
rect 197353 132502 200100 132504
rect 197353 132499 197419 132502
rect 369853 132426 369919 132429
rect 513465 132426 513531 132429
rect 369853 132424 369962 132426
rect 369853 132368 369858 132424
rect 369914 132368 369962 132424
rect 369853 132363 369962 132368
rect 171133 132290 171199 132293
rect 302509 132290 302575 132293
rect 169924 132288 171199 132290
rect 169924 132232 171138 132288
rect 171194 132232 171199 132288
rect 169924 132230 171199 132232
rect 299828 132288 302575 132290
rect 299828 132232 302514 132288
rect 302570 132232 302575 132288
rect 369902 132260 369962 132363
rect 513422 132424 513531 132426
rect 513422 132368 513470 132424
rect 513526 132368 513531 132424
rect 513422 132363 513531 132368
rect 513422 132260 513482 132363
rect 299828 132230 302575 132232
rect 171133 132227 171199 132230
rect 302509 132227 302575 132230
rect 444189 132154 444255 132157
rect 445109 132154 445175 132157
rect 441846 132152 445175 132154
rect 441846 132096 444194 132152
rect 444250 132096 445114 132152
rect 445170 132096 445175 132152
rect 441846 132094 445175 132096
rect 369485 132018 369551 132021
rect 369485 132016 369594 132018
rect 369485 131960 369490 132016
rect 369546 131960 369594 132016
rect 369485 131955 369594 131960
rect 172421 131746 172487 131749
rect 169924 131744 172487 131746
rect 169924 131688 172426 131744
rect 172482 131688 172487 131744
rect 369534 131716 369594 131955
rect 169924 131686 172487 131688
rect 172421 131683 172487 131686
rect 441846 131580 441906 132094
rect 444189 132091 444255 132094
rect 445109 132091 445175 132094
rect 514109 131746 514175 131749
rect 513820 131744 514175 131746
rect 513820 131688 514114 131744
rect 514170 131688 514175 131744
rect 513820 131686 514175 131688
rect 514109 131683 514175 131686
rect 369393 131474 369459 131477
rect 369350 131472 369459 131474
rect 369350 131416 369398 131472
rect 369454 131416 369459 131472
rect 369350 131411 369459 131416
rect 513557 131474 513623 131477
rect 513557 131472 513666 131474
rect 513557 131416 513562 131472
rect 513618 131416 513666 131472
rect 513557 131411 513666 131416
rect 172329 131202 172395 131205
rect 169924 131200 172395 131202
rect 169924 131144 172334 131200
rect 172390 131144 172395 131200
rect 369350 131172 369410 131411
rect 513606 131172 513666 131411
rect 169924 131142 172395 131144
rect 172329 131139 172395 131142
rect 171317 130658 171383 130661
rect 516133 130658 516199 130661
rect 169924 130656 171383 130658
rect 169924 130600 171322 130656
rect 171378 130600 171383 130656
rect 513820 130656 516199 130658
rect 169924 130598 171383 130600
rect 171317 130595 171383 130598
rect 197353 130386 197419 130389
rect 197353 130384 200100 130386
rect 197353 130328 197358 130384
rect 197414 130328 200100 130384
rect 197353 130326 200100 130328
rect 197353 130323 197419 130326
rect 369902 130250 369962 130628
rect 513820 130600 516138 130656
rect 516194 130600 516199 130656
rect 513820 130598 516199 130600
rect 516133 130595 516199 130598
rect 370037 130250 370103 130253
rect 369902 130248 370103 130250
rect 369902 130192 370042 130248
rect 370098 130192 370103 130248
rect 369902 130190 370103 130192
rect 370037 130187 370103 130190
rect 172237 130114 172303 130117
rect 370313 130114 370379 130117
rect 169924 130112 172303 130114
rect 169924 130056 172242 130112
rect 172298 130056 172303 130112
rect 169924 130054 172303 130056
rect 369932 130112 370379 130114
rect 369932 130056 370318 130112
rect 370374 130056 370379 130112
rect 369932 130054 370379 130056
rect 172237 130051 172303 130054
rect 370313 130051 370379 130054
rect 441846 129842 441906 130356
rect 516225 130114 516291 130117
rect 513820 130112 516291 130114
rect 513820 130056 516230 130112
rect 516286 130056 516291 130112
rect 513820 130054 516291 130056
rect 516225 130051 516291 130054
rect 442901 129842 442967 129845
rect 444465 129842 444531 129845
rect 441846 129840 444531 129842
rect 441846 129784 442906 129840
rect 442962 129784 444470 129840
rect 444526 129784 444531 129840
rect 441846 129782 444531 129784
rect 442901 129779 442967 129782
rect 444465 129779 444531 129782
rect 172421 129570 172487 129573
rect 373993 129570 374059 129573
rect 169924 129568 172487 129570
rect 169924 129512 172426 129568
rect 172482 129512 172487 129568
rect 369932 129568 374059 129570
rect 369932 129540 373998 129568
rect 169924 129510 172487 129512
rect 172421 129507 172487 129510
rect 369902 129512 373998 129540
rect 374054 129512 374059 129568
rect 369902 129510 374059 129512
rect 369902 129165 369962 129510
rect 373993 129507 374059 129510
rect 302693 129162 302759 129165
rect 299828 129160 302759 129162
rect 299828 129104 302698 129160
rect 302754 129104 302759 129160
rect 299828 129102 302759 129104
rect 302693 129099 302759 129102
rect 369853 129160 369962 129165
rect 369853 129104 369858 129160
rect 369914 129104 369962 129160
rect 369853 129102 369962 129104
rect 369853 129099 369919 129102
rect 172145 129026 172211 129029
rect 371785 129026 371851 129029
rect 169924 129024 172211 129026
rect 169924 128968 172150 129024
rect 172206 128968 172211 129024
rect 369380 129024 371851 129026
rect 369380 128996 371790 129024
rect 169924 128966 172211 128968
rect 172145 128963 172211 128966
rect 369350 128968 371790 128996
rect 371846 128968 371851 129024
rect 369350 128966 371851 128968
rect 369350 128621 369410 128966
rect 371785 128963 371851 128966
rect 441846 128754 441906 129268
rect 513281 129162 513347 129165
rect 513422 129162 513482 129540
rect 513281 129160 513482 129162
rect 513281 129104 513286 129160
rect 513342 129104 513482 129160
rect 513281 129102 513482 129104
rect 513281 129099 513347 129102
rect 443361 128754 443427 128757
rect 441846 128752 443427 128754
rect 441846 128696 443366 128752
rect 443422 128696 443427 128752
rect 441846 128694 443427 128696
rect 443361 128691 443427 128694
rect 513422 128621 513482 128996
rect 369301 128616 369410 128621
rect 369945 128618 370011 128621
rect 371877 128618 371943 128621
rect 369301 128560 369306 128616
rect 369362 128560 369410 128616
rect 369301 128558 369410 128560
rect 369902 128616 371943 128618
rect 369902 128560 369950 128616
rect 370006 128560 371882 128616
rect 371938 128560 371943 128616
rect 369902 128558 371943 128560
rect 513422 128616 513531 128621
rect 513422 128560 513470 128616
rect 513526 128560 513531 128616
rect 513422 128558 513531 128560
rect 369301 128555 369367 128558
rect 369902 128555 370011 128558
rect 371877 128555 371943 128558
rect 513465 128555 513531 128558
rect 171961 128482 172027 128485
rect 169924 128480 172027 128482
rect 169924 128424 171966 128480
rect 172022 128424 172027 128480
rect 369902 128452 369962 128555
rect 169924 128422 172027 128424
rect 171961 128419 172027 128422
rect 197353 128346 197419 128349
rect 197353 128344 200100 128346
rect 197353 128288 197358 128344
rect 197414 128288 200100 128344
rect 197353 128286 200100 128288
rect 197353 128283 197419 128286
rect 513790 128077 513850 128452
rect 444833 128074 444899 128077
rect 441876 128072 444899 128074
rect 441876 128044 444838 128072
rect 441846 128016 444838 128044
rect 444894 128016 444899 128072
rect 441846 128014 444899 128016
rect 513790 128072 513899 128077
rect 513790 128016 513838 128072
rect 513894 128016 513899 128072
rect 513790 128014 513899 128016
rect 172053 127938 172119 127941
rect 370221 127938 370287 127941
rect 372061 127938 372127 127941
rect 169924 127936 172119 127938
rect 169924 127880 172058 127936
rect 172114 127880 172119 127936
rect 169924 127878 172119 127880
rect 369932 127936 372127 127938
rect 369932 127880 370226 127936
rect 370282 127880 372066 127936
rect 372122 127880 372127 127936
rect 369932 127878 372127 127880
rect 172053 127875 172119 127878
rect 370221 127875 370287 127878
rect 372061 127875 372127 127878
rect 441846 127533 441906 128014
rect 444833 128011 444899 128014
rect 513833 128011 513899 128014
rect 513790 127533 513850 127908
rect 441846 127528 441955 127533
rect 441846 127472 441894 127528
rect 441950 127472 441955 127528
rect 441846 127470 441955 127472
rect 441889 127467 441955 127470
rect 513741 127528 513850 127533
rect 513741 127472 513746 127528
rect 513802 127472 513850 127528
rect 513741 127470 513850 127472
rect 513741 127467 513807 127470
rect 171777 127394 171843 127397
rect 370129 127394 370195 127397
rect 371918 127394 371924 127396
rect 169924 127392 171843 127394
rect 169924 127336 171782 127392
rect 171838 127336 171843 127392
rect 169924 127334 171843 127336
rect 369932 127392 371924 127394
rect 369932 127336 370134 127392
rect 370190 127336 371924 127392
rect 369932 127334 371924 127336
rect 171777 127331 171843 127334
rect 370129 127331 370195 127334
rect 371918 127332 371924 127334
rect 371988 127332 371994 127396
rect 513790 127122 513850 127364
rect 513925 127122 513991 127125
rect 513790 127120 513991 127122
rect 513790 127064 513930 127120
rect 513986 127064 513991 127120
rect 513790 127062 513991 127064
rect 513925 127059 513991 127062
rect 172329 126850 172395 126853
rect 169924 126848 172395 126850
rect 169924 126792 172334 126848
rect 172390 126792 172395 126848
rect 169924 126790 172395 126792
rect 172329 126787 172395 126790
rect 369350 126445 369410 126820
rect 441846 126445 441906 126956
rect 369350 126442 369459 126445
rect 371233 126442 371299 126445
rect 371693 126442 371759 126445
rect 369350 126440 371759 126442
rect 369350 126384 369398 126440
rect 369454 126384 371238 126440
rect 371294 126384 371698 126440
rect 371754 126384 371759 126440
rect 369350 126382 371759 126384
rect 369393 126379 369459 126382
rect 371233 126379 371299 126382
rect 371693 126379 371759 126382
rect 441797 126440 441906 126445
rect 441797 126384 441802 126440
rect 441858 126384 441906 126440
rect 441797 126382 441906 126384
rect 513790 126442 513850 126820
rect 514109 126442 514175 126445
rect 513790 126440 514175 126442
rect 513790 126384 514114 126440
rect 514170 126384 514175 126440
rect 513790 126382 514175 126384
rect 441797 126379 441863 126382
rect 514109 126379 514175 126382
rect 172421 126306 172487 126309
rect 370405 126306 370471 126309
rect 169924 126304 172487 126306
rect 169924 126248 172426 126304
rect 172482 126248 172487 126304
rect 169924 126246 172487 126248
rect 369932 126304 370471 126306
rect 369932 126248 370410 126304
rect 370466 126248 370471 126304
rect 369932 126246 370471 126248
rect 172421 126243 172487 126246
rect 370405 126243 370471 126246
rect 197629 126170 197695 126173
rect 302417 126170 302483 126173
rect 197629 126168 200100 126170
rect 197629 126112 197634 126168
rect 197690 126112 200100 126168
rect 197629 126110 200100 126112
rect 299828 126168 302483 126170
rect 299828 126112 302422 126168
rect 302478 126112 302483 126168
rect 299828 126110 302483 126112
rect 197629 126107 197695 126110
rect 302417 126107 302483 126110
rect 513606 125901 513666 126276
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 513606 125896 513715 125901
rect 513606 125840 513654 125896
rect 513710 125840 513715 125896
rect 583520 125884 584960 125974
rect 513606 125838 513715 125840
rect 513649 125835 513715 125838
rect 172237 125762 172303 125765
rect 370497 125762 370563 125765
rect 371601 125762 371667 125765
rect 442073 125762 442139 125765
rect 169924 125760 172303 125762
rect 169924 125704 172242 125760
rect 172298 125704 172303 125760
rect 169924 125702 172303 125704
rect 369932 125760 371667 125762
rect 369932 125704 370502 125760
rect 370558 125704 371606 125760
rect 371662 125704 371667 125760
rect 369932 125702 371667 125704
rect 441876 125760 442139 125762
rect 441876 125704 442078 125760
rect 442134 125704 442139 125760
rect 441876 125702 442139 125704
rect 172237 125699 172303 125702
rect 370497 125699 370563 125702
rect 371601 125699 371667 125702
rect 442073 125699 442139 125702
rect 513606 125357 513666 125732
rect 513373 125354 513439 125357
rect 513373 125352 513482 125354
rect 513373 125296 513378 125352
rect 513434 125296 513482 125352
rect 513373 125291 513482 125296
rect 513557 125352 513666 125357
rect 513557 125296 513562 125352
rect 513618 125296 513666 125352
rect 513557 125294 513666 125296
rect 513557 125291 513623 125294
rect 171501 125218 171567 125221
rect 371417 125218 371483 125221
rect 169924 125216 171567 125218
rect 169924 125160 171506 125216
rect 171562 125160 171567 125216
rect 169924 125158 171567 125160
rect 369932 125216 371483 125218
rect 369932 125160 371422 125216
rect 371478 125160 371483 125216
rect 513422 125188 513482 125291
rect 369932 125158 371483 125160
rect 171501 125155 171567 125158
rect 371417 125155 371483 125158
rect 441613 124946 441679 124949
rect 513373 124946 513439 124949
rect 441613 124944 441722 124946
rect 441613 124888 441618 124944
rect 441674 124888 441722 124944
rect 441613 124883 441722 124888
rect 513373 124944 513482 124946
rect 513373 124888 513378 124944
rect 513434 124888 513482 124944
rect 513373 124883 513482 124888
rect 171869 124674 171935 124677
rect 169924 124672 171935 124674
rect 169924 124616 171874 124672
rect 171930 124616 171935 124672
rect 441662 124644 441722 124883
rect 513422 124644 513482 124883
rect 169924 124614 171935 124616
rect 171869 124611 171935 124614
rect 369902 124405 369962 124644
rect 369853 124400 369962 124405
rect 369853 124344 369858 124400
rect 369914 124344 369962 124400
rect 369853 124342 369962 124344
rect 513281 124402 513347 124405
rect 513281 124400 513482 124402
rect 513281 124344 513286 124400
rect 513342 124344 513482 124400
rect 513281 124342 513482 124344
rect 369853 124339 369919 124342
rect 513281 124339 513347 124342
rect 172145 124266 172211 124269
rect 370865 124266 370931 124269
rect 169924 124264 172211 124266
rect 169924 124208 172150 124264
rect 172206 124208 172211 124264
rect 369932 124264 370931 124266
rect 369932 124236 370870 124264
rect 169924 124206 172211 124208
rect 172145 124203 172211 124206
rect 369902 124208 370870 124236
rect 370926 124208 370931 124264
rect 513422 124266 513482 124342
rect 517421 124266 517487 124269
rect 513422 124264 517487 124266
rect 513422 124236 517426 124264
rect 369902 124206 370931 124208
rect 513452 124208 517426 124236
rect 517482 124208 517487 124264
rect 513452 124206 517487 124208
rect 197353 124130 197419 124133
rect 197353 124128 200100 124130
rect 197353 124072 197358 124128
rect 197414 124072 200100 124128
rect 197353 124070 200100 124072
rect 197353 124067 197419 124070
rect 369902 123997 369962 124206
rect 370865 124203 370931 124206
rect 517421 124203 517487 124206
rect 362769 123996 362835 123997
rect 362718 123932 362724 123996
rect 362788 123994 362835 123996
rect 365161 123994 365227 123997
rect 365294 123994 365300 123996
rect 362788 123992 362880 123994
rect 362830 123936 362880 123992
rect 362788 123934 362880 123936
rect 365161 123992 365300 123994
rect 365161 123936 365166 123992
rect 365222 123936 365300 123992
rect 365161 123934 365300 123936
rect 362788 123932 362835 123934
rect 362769 123931 362835 123932
rect 365161 123931 365227 123934
rect 365294 123932 365300 123934
rect 365364 123932 365370 123996
rect 369902 123992 370011 123997
rect 369902 123936 369950 123992
rect 370006 123936 370011 123992
rect 369902 123934 370011 123936
rect 369945 123931 370011 123934
rect -960 123572 480 123812
rect 302233 123042 302299 123045
rect 299828 123040 302299 123042
rect 299828 122984 302238 123040
rect 302294 122984 302299 123040
rect 299828 122982 302299 122984
rect 302233 122979 302299 122982
rect 197445 121954 197511 121957
rect 197445 121952 200100 121954
rect 197445 121896 197450 121952
rect 197506 121896 200100 121952
rect 197445 121894 200100 121896
rect 197445 121891 197511 121894
rect 197353 119914 197419 119917
rect 302509 119914 302575 119917
rect 197353 119912 200100 119914
rect 197353 119856 197358 119912
rect 197414 119856 200100 119912
rect 197353 119854 200100 119856
rect 299828 119912 302575 119914
rect 299828 119856 302514 119912
rect 302570 119856 302575 119912
rect 299828 119854 302575 119856
rect 197353 119851 197419 119854
rect 302509 119851 302575 119854
rect 197629 117738 197695 117741
rect 197629 117736 200100 117738
rect 197629 117680 197634 117736
rect 197690 117680 200100 117736
rect 197629 117678 200100 117680
rect 197629 117675 197695 117678
rect 302601 116922 302667 116925
rect 299828 116920 302667 116922
rect 299828 116864 302606 116920
rect 302662 116864 302667 116920
rect 299828 116862 302667 116864
rect 302601 116859 302667 116862
rect 198549 115698 198615 115701
rect 198549 115696 200100 115698
rect 198549 115640 198554 115696
rect 198610 115640 200100 115696
rect 198549 115638 200100 115640
rect 198549 115635 198615 115638
rect 302969 113794 303035 113797
rect 299828 113792 303035 113794
rect 299828 113736 302974 113792
rect 303030 113736 303035 113792
rect 299828 113734 303035 113736
rect 302969 113731 303035 113734
rect 197537 113522 197603 113525
rect 197537 113520 200100 113522
rect 197537 113464 197542 113520
rect 197598 113464 200100 113520
rect 197537 113462 200100 113464
rect 197537 113459 197603 113462
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 197353 111482 197419 111485
rect 197353 111480 200100 111482
rect 197353 111424 197358 111480
rect 197414 111424 200100 111480
rect 197353 111422 200100 111424
rect 197353 111419 197419 111422
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect 302509 110666 302575 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect 299828 110664 302575 110666
rect 299828 110608 302514 110664
rect 302570 110608 302575 110664
rect 299828 110606 302575 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 302509 110603 302575 110606
rect 197537 109306 197603 109309
rect 197537 109304 200100 109306
rect 197537 109248 197542 109304
rect 197598 109248 200100 109304
rect 197537 109246 200100 109248
rect 197537 109243 197603 109246
rect 302785 107674 302851 107677
rect 299828 107672 302851 107674
rect 299828 107616 302790 107672
rect 302846 107616 302851 107672
rect 299828 107614 302851 107616
rect 302785 107611 302851 107614
rect 197997 107266 198063 107269
rect 197997 107264 200100 107266
rect 197997 107208 198002 107264
rect 198058 107208 200100 107264
rect 197997 107206 200100 107208
rect 197997 107203 198063 107206
rect 197445 105090 197511 105093
rect 197445 105088 200100 105090
rect 197445 105032 197450 105088
rect 197506 105032 200100 105088
rect 197445 105030 200100 105032
rect 197445 105027 197511 105030
rect 302877 104546 302943 104549
rect 299828 104544 302943 104546
rect 299828 104488 302882 104544
rect 302938 104488 302943 104544
rect 299828 104486 302943 104488
rect 302877 104483 302943 104486
rect 197997 103050 198063 103053
rect 197997 103048 200100 103050
rect 197997 102992 198002 103048
rect 198058 102992 200100 103048
rect 197997 102990 200100 102992
rect 197997 102987 198063 102990
rect 302785 101554 302851 101557
rect 299828 101552 302851 101554
rect 299828 101496 302790 101552
rect 302846 101496 302851 101552
rect 299828 101494 302851 101496
rect 302785 101491 302851 101494
rect 197997 101010 198063 101013
rect 197997 101008 200100 101010
rect 197997 100952 198002 101008
rect 198058 100952 200100 101008
rect 197997 100950 200100 100952
rect 197997 100947 198063 100950
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 195329 97882 195395 97885
rect 200849 97882 200915 97885
rect 195329 97880 200915 97882
rect 195329 97824 195334 97880
rect 195390 97824 200854 97880
rect 200910 97824 200915 97880
rect 195329 97822 200915 97824
rect 195329 97819 195395 97822
rect 200849 97819 200915 97822
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 281993 97610 282059 97613
rect 285857 97610 285923 97613
rect 281993 97608 285923 97610
rect 281993 97552 281998 97608
rect 282054 97552 285862 97608
rect 285918 97552 285923 97608
rect 281993 97550 285923 97552
rect 281993 97547 282059 97550
rect 285857 97547 285923 97550
rect 297909 97474 297975 97477
rect 450537 97474 450603 97477
rect 297909 97472 450603 97474
rect 297909 97416 297914 97472
rect 297970 97416 450542 97472
rect 450598 97416 450603 97472
rect 297909 97414 450603 97416
rect 297909 97411 297975 97414
rect 450537 97411 450603 97414
rect 280153 97338 280219 97341
rect 447777 97338 447843 97341
rect 280153 97336 447843 97338
rect 280153 97280 280158 97336
rect 280214 97280 447782 97336
rect 447838 97280 447843 97336
rect 280153 97278 447843 97280
rect 280153 97275 280219 97278
rect 447777 97275 447843 97278
rect 39297 97202 39363 97205
rect 203425 97202 203491 97205
rect 39297 97200 203491 97202
rect 39297 97144 39302 97200
rect 39358 97144 203430 97200
rect 203486 97144 203491 97200
rect 39297 97142 203491 97144
rect 39297 97139 39363 97142
rect 203425 97139 203491 97142
rect 297725 97202 297791 97205
rect 580257 97202 580323 97205
rect 297725 97200 580323 97202
rect 297725 97144 297730 97200
rect 297786 97144 580262 97200
rect 580318 97144 580323 97200
rect 297725 97142 580323 97144
rect 297725 97139 297791 97142
rect 580257 97139 580323 97142
rect 297081 96658 297147 96661
rect 298737 96658 298803 96661
rect 297081 96656 298803 96658
rect 297081 96600 297086 96656
rect 297142 96600 298742 96656
rect 298798 96600 298803 96656
rect 297081 96598 298803 96600
rect 297081 96595 297147 96598
rect 298737 96595 298803 96598
rect 289905 95978 289971 95981
rect 532693 95978 532759 95981
rect 289905 95976 532759 95978
rect 289905 95920 289910 95976
rect 289966 95920 532698 95976
rect 532754 95920 532759 95976
rect 289905 95918 532759 95920
rect 289905 95915 289971 95918
rect 532693 95915 532759 95918
rect 293125 95842 293191 95845
rect 547137 95842 547203 95845
rect 293125 95840 547203 95842
rect 293125 95784 293130 95840
rect 293186 95784 547142 95840
rect 547198 95784 547203 95840
rect 293125 95782 547203 95784
rect 293125 95779 293191 95782
rect 547137 95779 547203 95782
rect 12341 94482 12407 94485
rect 202045 94482 202111 94485
rect 12341 94480 202111 94482
rect 12341 94424 12346 94480
rect 12402 94424 202050 94480
rect 202106 94424 202111 94480
rect 12341 94422 202111 94424
rect 12341 94419 12407 94422
rect 202045 94419 202111 94422
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 582465 46338 582531 46341
rect 583520 46338 584960 46428
rect 582465 46336 584960 46338
rect 582465 46280 582470 46336
rect 582526 46280 584960 46336
rect 582465 46278 584960 46280
rect 582465 46275 582531 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 371188 584020 371252 584084
rect 371372 583476 371436 583540
rect 371556 582932 371620 582996
rect 371740 572188 371804 572252
rect 361620 553420 361684 553484
rect 365300 553420 365364 553484
rect 435220 553480 435284 553484
rect 435220 553424 435234 553480
rect 435234 553424 435284 553480
rect 435220 553420 435284 553424
rect 436692 553480 436756 553484
rect 436692 553424 436742 553480
rect 436742 553424 436756 553480
rect 436692 553420 436756 553424
rect 444604 511532 444668 511596
rect 444788 500788 444852 500852
rect 444420 500244 444484 500308
rect 365300 484060 365364 484124
rect 435220 483984 435284 483988
rect 435220 483928 435234 483984
rect 435234 483928 435284 483984
rect 435220 483924 435284 483928
rect 436692 483984 436756 483988
rect 436692 483928 436742 483984
rect 436742 483928 436756 483984
rect 436692 483924 436756 483928
rect 365300 482836 365364 482900
rect 361620 482156 361684 482220
rect 362724 482156 362788 482220
rect 371188 439996 371252 440060
rect 371372 439452 371436 439516
rect 516180 439452 516244 439516
rect 371188 439044 371252 439108
rect 372476 439044 372540 439108
rect 371188 438908 371252 438972
rect 371556 438908 371620 438972
rect 371924 428708 371988 428772
rect 371740 428164 371804 428228
rect 369348 427348 369412 427412
rect 362724 412040 362788 412044
rect 362724 411984 362774 412040
rect 362774 411984 362788 412040
rect 362724 411980 362788 411984
rect 365300 411980 365364 412044
rect 440740 409532 440804 409596
rect 361620 409124 361684 409188
rect 362724 409124 362788 409188
rect 434852 408640 434916 408644
rect 434852 408584 434902 408640
rect 434902 408584 434916 408640
rect 434852 408580 434916 408584
rect 436140 408580 436204 408644
rect 444604 367508 444668 367572
rect 444420 357172 444484 357236
rect 444604 356764 444668 356828
rect 444420 356220 444484 356284
rect 444788 354588 444852 354652
rect 361620 340444 361684 340508
rect 364380 340444 364444 340508
rect 366588 340444 366652 340508
rect 436140 340036 436204 340100
rect 440740 340096 440804 340100
rect 440740 340040 440790 340096
rect 440790 340040 440804 340096
rect 440740 340036 440804 340040
rect 434852 339960 434916 339964
rect 434852 339904 434856 339960
rect 434856 339904 434912 339960
rect 434912 339904 434916 339960
rect 434852 339900 434916 339904
rect 216812 299372 216876 299436
rect 216812 299100 216876 299164
rect 516364 298148 516428 298212
rect 371372 298012 371436 298076
rect 371924 298012 371988 298076
rect 372476 296108 372540 296172
rect 516180 295836 516244 295900
rect 371556 295292 371620 295356
rect 371740 295292 371804 295356
rect 371188 295020 371252 295084
rect 516364 293796 516428 293860
rect 372292 289852 372356 289916
rect 372108 289444 372172 289508
rect 369348 283868 369412 283932
rect 371924 269860 371988 269924
rect 444604 267684 444668 267748
rect 361620 266188 361684 266252
rect 364380 265780 364444 265844
rect 436692 265508 436756 265572
rect 435220 264964 435284 265028
rect 372292 231780 372356 231844
rect 372108 231644 372172 231708
rect 365116 225660 365180 225724
rect 366588 225660 366652 225724
rect 444604 212740 444668 212804
rect 444788 212332 444852 212396
rect 444420 212196 444484 212260
rect 444788 211108 444852 211172
rect 371924 203492 371988 203556
rect 444420 201180 444484 201244
rect 444604 198868 444668 198932
rect 365300 196420 365364 196484
rect 366588 196420 366652 196484
rect 435220 196072 435284 196076
rect 435220 196016 435234 196072
rect 435234 196016 435284 196072
rect 435220 196012 435284 196016
rect 436692 196072 436756 196076
rect 436692 196016 436742 196072
rect 436742 196016 436756 196072
rect 436692 196012 436756 196016
rect 361620 194516 361684 194580
rect 362724 194516 362788 194580
rect 444788 169628 444852 169692
rect 444788 168948 444852 169012
rect 371924 158748 371988 158812
rect 444604 158748 444668 158812
rect 444788 156436 444852 156500
rect 372108 153716 372172 153780
rect 372292 153172 372356 153236
rect 371188 152960 371252 152964
rect 371188 152904 371238 152960
rect 371238 152904 371252 152960
rect 371188 152900 371252 152904
rect 514156 152900 514220 152964
rect 371556 152628 371620 152692
rect 371740 152084 371804 152148
rect 513972 152356 514036 152420
rect 514340 152008 514404 152012
rect 514340 151952 514390 152008
rect 514390 151952 514404 152008
rect 514340 151948 514404 151952
rect 514156 151812 514220 151876
rect 514340 151404 514404 151468
rect 513972 151268 514036 151332
rect 371188 148276 371252 148340
rect 444420 134948 444484 135012
rect 371924 127332 371988 127396
rect 362724 123992 362788 123996
rect 362724 123936 362774 123992
rect 362774 123936 362788 123992
rect 362724 123932 362788 123936
rect 365300 123932 365364 123996
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 192000 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 192000 168134 204618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 192000 171854 208338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 162243 183454 162563 183486
rect 162243 183218 162285 183454
rect 162521 183218 162563 183454
rect 162243 183134 162563 183218
rect 162243 182898 162285 183134
rect 162521 182898 162563 183134
rect 162243 182866 162563 182898
rect 164840 183454 165160 183486
rect 164840 183218 164882 183454
rect 165118 183218 165160 183454
rect 164840 183134 165160 183218
rect 164840 182898 164882 183134
rect 165118 182898 165160 183134
rect 164840 182866 165160 182898
rect 167437 183454 167757 183486
rect 167437 183218 167479 183454
rect 167715 183218 167757 183454
rect 167437 183134 167757 183218
rect 167437 182898 167479 183134
rect 167715 182898 167757 183134
rect 167437 182866 167757 182898
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 163541 165454 163861 165486
rect 163541 165218 163583 165454
rect 163819 165218 163861 165454
rect 163541 165134 163861 165218
rect 163541 164898 163583 165134
rect 163819 164898 163861 165134
rect 163541 164866 163861 164898
rect 166138 165454 166458 165486
rect 166138 165218 166180 165454
rect 166416 165218 166458 165454
rect 166138 165134 166458 165218
rect 166138 164898 166180 165134
rect 166416 164898 166458 165134
rect 166138 164866 166458 164898
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 163794 156000 164414 158000
rect 167514 156000 168134 158000
rect 171234 156000 171854 158000
rect 162243 147454 162563 147486
rect 162243 147218 162285 147454
rect 162521 147218 162563 147454
rect 162243 147134 162563 147218
rect 162243 146898 162285 147134
rect 162521 146898 162563 147134
rect 162243 146866 162563 146898
rect 164840 147454 165160 147486
rect 164840 147218 164882 147454
rect 165118 147218 165160 147454
rect 164840 147134 165160 147218
rect 164840 146898 164882 147134
rect 165118 146898 165160 147134
rect 164840 146866 165160 146898
rect 167437 147454 167757 147486
rect 167437 147218 167479 147454
rect 167715 147218 167757 147454
rect 167437 147134 167757 147218
rect 167437 146898 167479 147134
rect 167715 146898 167757 147134
rect 167437 146866 167757 146898
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 163541 129454 163861 129486
rect 163541 129218 163583 129454
rect 163819 129218 163861 129454
rect 163541 129134 163861 129218
rect 163541 128898 163583 129134
rect 163819 128898 163861 129134
rect 163541 128866 163861 128898
rect 166138 129454 166458 129486
rect 166138 129218 166180 129454
rect 166416 129218 166458 129454
rect 166138 129134 166458 129218
rect 166138 128898 166180 129134
rect 166416 128898 166458 129134
rect 166138 128866 166458 128898
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 93454 164414 122000
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 97174 168134 122000
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 100894 171854 122000
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 302000 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 302000 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 302000 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 302000 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 302000 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 302000 222134 330618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 302000 225854 334338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 302000 229574 302058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 302000 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 302000 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 302000 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 302000 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 302000 254414 326898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 302000 258134 330618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 302000 261854 334338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 302000 265574 302058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 302000 272414 308898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 302000 276134 312618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 302000 279854 316338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 302000 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 302000 290414 326898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 302000 294134 330618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 302000 297854 334338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 302000 301574 302058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 216811 299436 216877 299437
rect 216811 299372 216812 299436
rect 216876 299372 216877 299436
rect 216811 299371 216877 299372
rect 216814 299165 216874 299371
rect 216811 299164 216877 299165
rect 216811 299100 216812 299164
rect 216876 299100 216877 299164
rect 216811 299099 216877 299100
rect 204208 291454 204528 291486
rect 204208 291218 204250 291454
rect 204486 291218 204528 291454
rect 204208 291134 204528 291218
rect 204208 290898 204250 291134
rect 204486 290898 204528 291134
rect 204208 290866 204528 290898
rect 234928 291454 235248 291486
rect 234928 291218 234970 291454
rect 235206 291218 235248 291454
rect 234928 291134 235248 291218
rect 234928 290898 234970 291134
rect 235206 290898 235248 291134
rect 234928 290866 235248 290898
rect 265648 291454 265968 291486
rect 265648 291218 265690 291454
rect 265926 291218 265968 291454
rect 265648 291134 265968 291218
rect 265648 290898 265690 291134
rect 265926 290898 265968 291134
rect 265648 290866 265968 290898
rect 296368 291454 296688 291486
rect 296368 291218 296410 291454
rect 296646 291218 296688 291454
rect 296368 291134 296688 291218
rect 296368 290898 296410 291134
rect 296646 290898 296688 291134
rect 296368 290866 296688 290898
rect 219568 273454 219888 273486
rect 219568 273218 219610 273454
rect 219846 273218 219888 273454
rect 219568 273134 219888 273218
rect 219568 272898 219610 273134
rect 219846 272898 219888 273134
rect 219568 272866 219888 272898
rect 250288 273454 250608 273486
rect 250288 273218 250330 273454
rect 250566 273218 250608 273454
rect 250288 273134 250608 273218
rect 250288 272898 250330 273134
rect 250566 272898 250608 273134
rect 250288 272866 250608 272898
rect 281008 273454 281328 273486
rect 281008 273218 281050 273454
rect 281286 273218 281328 273454
rect 281008 273134 281328 273218
rect 281008 272898 281050 273134
rect 281286 272898 281328 273134
rect 281008 272866 281328 272898
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 204208 255454 204528 255486
rect 204208 255218 204250 255454
rect 204486 255218 204528 255454
rect 204208 255134 204528 255218
rect 204208 254898 204250 255134
rect 204486 254898 204528 255134
rect 204208 254866 204528 254898
rect 234928 255454 235248 255486
rect 234928 255218 234970 255454
rect 235206 255218 235248 255454
rect 234928 255134 235248 255218
rect 234928 254898 234970 255134
rect 235206 254898 235248 255134
rect 234928 254866 235248 254898
rect 265648 255454 265968 255486
rect 265648 255218 265690 255454
rect 265926 255218 265968 255454
rect 265648 255134 265968 255218
rect 265648 254898 265690 255134
rect 265926 254898 265968 255134
rect 265648 254866 265968 254898
rect 296368 255454 296688 255486
rect 296368 255218 296410 255454
rect 296646 255218 296688 255454
rect 296368 255134 296688 255218
rect 296368 254898 296410 255134
rect 296646 254898 296688 255134
rect 296368 254866 296688 254898
rect 219568 237454 219888 237486
rect 219568 237218 219610 237454
rect 219846 237218 219888 237454
rect 219568 237134 219888 237218
rect 219568 236898 219610 237134
rect 219846 236898 219888 237134
rect 219568 236866 219888 236898
rect 250288 237454 250608 237486
rect 250288 237218 250330 237454
rect 250566 237218 250608 237454
rect 250288 237134 250608 237218
rect 250288 236898 250330 237134
rect 250566 236898 250608 237134
rect 250288 236866 250608 236898
rect 281008 237454 281328 237486
rect 281008 237218 281050 237454
rect 281286 237218 281328 237454
rect 281008 237134 281328 237218
rect 281008 236898 281050 237134
rect 281286 236898 281328 237134
rect 281008 236866 281328 236898
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 204208 219454 204528 219486
rect 204208 219218 204250 219454
rect 204486 219218 204528 219454
rect 204208 219134 204528 219218
rect 204208 218898 204250 219134
rect 204486 218898 204528 219134
rect 204208 218866 204528 218898
rect 234928 219454 235248 219486
rect 234928 219218 234970 219454
rect 235206 219218 235248 219454
rect 234928 219134 235248 219218
rect 234928 218898 234970 219134
rect 235206 218898 235248 219134
rect 234928 218866 235248 218898
rect 265648 219454 265968 219486
rect 265648 219218 265690 219454
rect 265926 219218 265968 219454
rect 265648 219134 265968 219218
rect 265648 218898 265690 219134
rect 265926 218898 265968 219134
rect 265648 218866 265968 218898
rect 296368 219454 296688 219486
rect 296368 219218 296410 219454
rect 296646 219218 296688 219454
rect 296368 219134 296688 219218
rect 296368 218898 296410 219134
rect 296646 218898 296688 219134
rect 296368 218866 296688 218898
rect 219568 201454 219888 201486
rect 219568 201218 219610 201454
rect 219846 201218 219888 201454
rect 219568 201134 219888 201218
rect 219568 200898 219610 201134
rect 219846 200898 219888 201134
rect 219568 200866 219888 200898
rect 250288 201454 250608 201486
rect 250288 201218 250330 201454
rect 250566 201218 250608 201454
rect 250288 201134 250608 201218
rect 250288 200898 250330 201134
rect 250566 200898 250608 201134
rect 250288 200866 250608 200898
rect 281008 201454 281328 201486
rect 281008 201218 281050 201454
rect 281286 201218 281328 201454
rect 281008 201134 281328 201218
rect 281008 200898 281050 201134
rect 281286 200898 281328 201134
rect 281008 200866 281328 200898
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 204208 183454 204528 183486
rect 204208 183218 204250 183454
rect 204486 183218 204528 183454
rect 204208 183134 204528 183218
rect 204208 182898 204250 183134
rect 204486 182898 204528 183134
rect 204208 182866 204528 182898
rect 234928 183454 235248 183486
rect 234928 183218 234970 183454
rect 235206 183218 235248 183454
rect 234928 183134 235248 183218
rect 234928 182898 234970 183134
rect 235206 182898 235248 183134
rect 234928 182866 235248 182898
rect 265648 183454 265968 183486
rect 265648 183218 265690 183454
rect 265926 183218 265968 183454
rect 265648 183134 265968 183218
rect 265648 182898 265690 183134
rect 265926 182898 265968 183134
rect 265648 182866 265968 182898
rect 296368 183454 296688 183486
rect 296368 183218 296410 183454
rect 296646 183218 296688 183454
rect 296368 183134 296688 183218
rect 296368 182898 296410 183134
rect 296646 182898 296688 183134
rect 296368 182866 296688 182898
rect 219568 165454 219888 165486
rect 219568 165218 219610 165454
rect 219846 165218 219888 165454
rect 219568 165134 219888 165218
rect 219568 164898 219610 165134
rect 219846 164898 219888 165134
rect 219568 164866 219888 164898
rect 250288 165454 250608 165486
rect 250288 165218 250330 165454
rect 250566 165218 250608 165454
rect 250288 165134 250608 165218
rect 250288 164898 250330 165134
rect 250566 164898 250608 165134
rect 250288 164866 250608 164898
rect 281008 165454 281328 165486
rect 281008 165218 281050 165454
rect 281286 165218 281328 165454
rect 281008 165134 281328 165218
rect 281008 164898 281050 165134
rect 281286 164898 281328 165134
rect 281008 164866 281328 164898
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 204208 147454 204528 147486
rect 204208 147218 204250 147454
rect 204486 147218 204528 147454
rect 204208 147134 204528 147218
rect 204208 146898 204250 147134
rect 204486 146898 204528 147134
rect 204208 146866 204528 146898
rect 234928 147454 235248 147486
rect 234928 147218 234970 147454
rect 235206 147218 235248 147454
rect 234928 147134 235248 147218
rect 234928 146898 234970 147134
rect 235206 146898 235248 147134
rect 234928 146866 235248 146898
rect 265648 147454 265968 147486
rect 265648 147218 265690 147454
rect 265926 147218 265968 147454
rect 265648 147134 265968 147218
rect 265648 146898 265690 147134
rect 265926 146898 265968 147134
rect 265648 146866 265968 146898
rect 296368 147454 296688 147486
rect 296368 147218 296410 147454
rect 296646 147218 296688 147454
rect 296368 147134 296688 147218
rect 296368 146898 296410 147134
rect 296646 146898 296688 147134
rect 296368 146866 296688 146898
rect 219568 129454 219888 129486
rect 219568 129218 219610 129454
rect 219846 129218 219888 129454
rect 219568 129134 219888 129218
rect 219568 128898 219610 129134
rect 219846 128898 219888 129134
rect 219568 128866 219888 128898
rect 250288 129454 250608 129486
rect 250288 129218 250330 129454
rect 250566 129218 250608 129454
rect 250288 129134 250608 129218
rect 250288 128898 250330 129134
rect 250566 128898 250608 129134
rect 250288 128866 250608 128898
rect 281008 129454 281328 129486
rect 281008 129218 281050 129454
rect 281286 129218 281328 129454
rect 281008 129134 281328 129218
rect 281008 128898 281050 129134
rect 281286 128898 281328 129134
rect 281008 128866 281328 128898
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 204208 111454 204528 111486
rect 204208 111218 204250 111454
rect 204486 111218 204528 111454
rect 204208 111134 204528 111218
rect 204208 110898 204250 111134
rect 204486 110898 204528 111134
rect 204208 110866 204528 110898
rect 234928 111454 235248 111486
rect 234928 111218 234970 111454
rect 235206 111218 235248 111454
rect 234928 111134 235248 111218
rect 234928 110898 234970 111134
rect 235206 110898 235248 111134
rect 234928 110866 235248 110898
rect 265648 111454 265968 111486
rect 265648 111218 265690 111454
rect 265926 111218 265968 111454
rect 265648 111134 265968 111218
rect 265648 110898 265690 111134
rect 265926 110898 265968 111134
rect 265648 110866 265968 110898
rect 296368 111454 296688 111486
rect 296368 111218 296410 111454
rect 296646 111218 296688 111454
rect 296368 111134 296688 111218
rect 296368 110898 296410 111134
rect 296646 110898 296688 111134
rect 296368 110866 296688 110898
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 98000
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 97174 204134 98000
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 98000
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 98000
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 98000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 98000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 98000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 98000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 98000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 98000
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 98000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 98000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 98000
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 98000
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 82894 261854 98000
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 86614 265574 98000
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 98000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 97174 276134 98000
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 98000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 98000
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 98000
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 79174 294134 98000
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 98000
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 86614 301574 98000
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 588000 362414 614898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 588000 366134 618618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 588000 369854 622338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 371187 584084 371253 584085
rect 371187 584020 371188 584084
rect 371252 584020 371253 584084
rect 371187 584019 371253 584020
rect 362243 579454 362563 579486
rect 362243 579218 362285 579454
rect 362521 579218 362563 579454
rect 362243 579134 362563 579218
rect 362243 578898 362285 579134
rect 362521 578898 362563 579134
rect 362243 578866 362563 578898
rect 364840 579454 365160 579486
rect 364840 579218 364882 579454
rect 365118 579218 365160 579454
rect 364840 579134 365160 579218
rect 364840 578898 364882 579134
rect 365118 578898 365160 579134
rect 364840 578866 365160 578898
rect 367437 579454 367757 579486
rect 367437 579218 367479 579454
rect 367715 579218 367757 579454
rect 367437 579134 367757 579218
rect 367437 578898 367479 579134
rect 367715 578898 367757 579134
rect 367437 578866 367757 578898
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 363541 561454 363861 561486
rect 363541 561218 363583 561454
rect 363819 561218 363861 561454
rect 363541 561134 363861 561218
rect 363541 560898 363583 561134
rect 363819 560898 363861 561134
rect 363541 560866 363861 560898
rect 366138 561454 366458 561486
rect 366138 561218 366180 561454
rect 366416 561218 366458 561454
rect 366138 561134 366458 561218
rect 366138 560898 366180 561134
rect 366416 560898 366458 561134
rect 366138 560866 366458 560898
rect 361619 553484 361685 553485
rect 361619 553420 361620 553484
rect 361684 553420 361685 553484
rect 361619 553419 361685 553420
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 361622 482221 361682 553419
rect 361794 543454 362414 554000
rect 365299 553484 365365 553485
rect 365299 553420 365300 553484
rect 365364 553420 365365 553484
rect 365299 553419 365365 553420
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 516000 362414 542898
rect 365302 520290 365362 553419
rect 365118 520230 365362 520290
rect 365514 547174 366134 554000
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365118 512010 365178 520230
rect 365514 516000 366134 546618
rect 369234 550894 369854 554000
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 516000 369854 550338
rect 365118 511950 366650 512010
rect 362243 507454 362563 507486
rect 362243 507218 362285 507454
rect 362521 507218 362563 507454
rect 362243 507134 362563 507218
rect 362243 506898 362285 507134
rect 362521 506898 362563 507134
rect 362243 506866 362563 506898
rect 364840 507454 365160 507486
rect 364840 507218 364882 507454
rect 365118 507218 365160 507454
rect 364840 507134 365160 507218
rect 364840 506898 364882 507134
rect 365118 506898 365160 507134
rect 364840 506866 365160 506898
rect 363541 489454 363861 489486
rect 363541 489218 363583 489454
rect 363819 489218 363861 489454
rect 363541 489134 363861 489218
rect 363541 488898 363583 489134
rect 363819 488898 363861 489134
rect 363541 488866 363861 488898
rect 366138 489454 366458 489486
rect 366138 489218 366180 489454
rect 366416 489218 366458 489454
rect 366138 489134 366458 489218
rect 366138 488898 366180 489134
rect 366416 488898 366458 489134
rect 366138 488866 366458 488898
rect 366590 485790 366650 511950
rect 367437 507454 367757 507486
rect 367437 507218 367479 507454
rect 367715 507218 367757 507454
rect 367437 507134 367757 507218
rect 367437 506898 367479 507134
rect 367715 506898 367757 507134
rect 367437 506866 367757 506898
rect 365118 485730 366650 485790
rect 365118 484394 365178 485730
rect 365118 484334 365362 484394
rect 365302 484125 365362 484334
rect 365299 484124 365365 484125
rect 365299 484060 365300 484124
rect 365364 484060 365365 484124
rect 365299 484059 365365 484060
rect 365302 482901 365362 484059
rect 365299 482900 365365 482901
rect 365299 482836 365300 482900
rect 365364 482836 365365 482900
rect 365299 482835 365365 482836
rect 361619 482220 361685 482221
rect 361619 482156 361620 482220
rect 361684 482156 361685 482220
rect 361619 482155 361685 482156
rect 362723 482220 362789 482221
rect 362723 482156 362724 482220
rect 362788 482156 362789 482220
rect 362723 482155 362789 482156
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 361794 471454 362414 482000
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 444000 362414 470898
rect 362243 435454 362563 435486
rect 362243 435218 362285 435454
rect 362521 435218 362563 435454
rect 362243 435134 362563 435218
rect 362243 434898 362285 435134
rect 362521 434898 362563 435134
rect 362243 434866 362563 434898
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 362726 412045 362786 482155
rect 364840 435454 365160 435486
rect 364840 435218 364882 435454
rect 365118 435218 365160 435454
rect 364840 435134 365160 435218
rect 364840 434898 364882 435134
rect 365118 434898 365160 435134
rect 364840 434866 365160 434898
rect 363541 417454 363861 417486
rect 363541 417218 363583 417454
rect 363819 417218 363861 417454
rect 363541 417134 363861 417218
rect 363541 416898 363583 417134
rect 363819 416898 363861 417134
rect 363541 416866 363861 416898
rect 365302 412045 365362 482835
rect 365514 475174 366134 482000
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 444000 366134 474618
rect 369234 478894 369854 482000
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 444000 369854 478338
rect 371190 440061 371250 584019
rect 371371 583540 371437 583541
rect 371371 583476 371372 583540
rect 371436 583476 371437 583540
rect 371371 583475 371437 583476
rect 371187 440060 371253 440061
rect 371187 439996 371188 440060
rect 371252 439996 371253 440060
rect 371187 439995 371253 439996
rect 371190 439109 371250 439995
rect 371374 439517 371434 583475
rect 371555 582996 371621 582997
rect 371555 582932 371556 582996
rect 371620 582932 371621 582996
rect 371555 582931 371621 582932
rect 371371 439516 371437 439517
rect 371371 439452 371372 439516
rect 371436 439452 371437 439516
rect 371371 439451 371437 439452
rect 371187 439108 371253 439109
rect 371187 439044 371188 439108
rect 371252 439044 371253 439108
rect 371187 439043 371253 439044
rect 371187 438972 371253 438973
rect 371187 438908 371188 438972
rect 371252 438908 371253 438972
rect 371187 438907 371253 438908
rect 367437 435454 367757 435486
rect 367437 435218 367479 435454
rect 367715 435218 367757 435454
rect 367437 435134 367757 435218
rect 367437 434898 367479 435134
rect 367715 434898 367757 435134
rect 367437 434866 367757 434898
rect 369347 427412 369413 427413
rect 369347 427348 369348 427412
rect 369412 427348 369413 427412
rect 369347 427347 369413 427348
rect 366138 417454 366458 417486
rect 366138 417218 366180 417454
rect 366416 417218 366458 417454
rect 366138 417134 366458 417218
rect 366138 416898 366180 417134
rect 366416 416898 366458 417134
rect 366138 416866 366458 416898
rect 369350 412650 369410 427347
rect 368430 412590 369410 412650
rect 362723 412044 362789 412045
rect 362723 411980 362724 412044
rect 362788 411980 362789 412044
rect 362723 411979 362789 411980
rect 365299 412044 365365 412045
rect 365299 411980 365300 412044
rect 365364 411980 365365 412044
rect 365299 411979 365365 411980
rect 361619 409188 361685 409189
rect 361619 409124 361620 409188
rect 361684 409124 361685 409188
rect 361619 409123 361685 409124
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 361622 340509 361682 409123
rect 361794 399454 362414 410000
rect 362726 409189 362786 411979
rect 362723 409188 362789 409189
rect 362723 409124 362724 409188
rect 362788 409124 362789 409188
rect 362723 409123 362789 409124
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 372000 362414 398898
rect 365302 376770 365362 411979
rect 364750 376710 365362 376770
rect 365514 403174 366134 410000
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 364750 368490 364810 376710
rect 365514 372000 366134 402618
rect 368430 368490 368490 412590
rect 369234 406894 369854 410000
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 372000 369854 406338
rect 364750 368430 366650 368490
rect 362243 363454 362563 363486
rect 362243 363218 362285 363454
rect 362521 363218 362563 363454
rect 362243 363134 362563 363218
rect 362243 362898 362285 363134
rect 362521 362898 362563 363134
rect 362243 362866 362563 362898
rect 364840 363454 365160 363486
rect 364840 363218 364882 363454
rect 365118 363218 365160 363454
rect 364840 363134 365160 363218
rect 364840 362898 364882 363134
rect 365118 362898 365160 363134
rect 364840 362866 365160 362898
rect 363541 345454 363861 345486
rect 363541 345218 363583 345454
rect 363819 345218 363861 345454
rect 363541 345134 363861 345218
rect 363541 344898 363583 345134
rect 363819 344898 363861 345134
rect 363541 344866 363861 344898
rect 366138 345454 366458 345486
rect 366138 345218 366180 345454
rect 366416 345218 366458 345454
rect 366138 345134 366458 345218
rect 366138 344898 366180 345134
rect 366416 344898 366458 345134
rect 366138 344866 366458 344898
rect 366590 340509 366650 368430
rect 368246 368430 368490 368490
rect 367437 363454 367757 363486
rect 367437 363218 367479 363454
rect 367715 363218 367757 363454
rect 367437 363134 367757 363218
rect 367437 362898 367479 363134
rect 367715 362898 367757 363134
rect 367437 362866 367757 362898
rect 361619 340508 361685 340509
rect 361619 340444 361620 340508
rect 361684 340444 361685 340508
rect 361619 340443 361685 340444
rect 364379 340508 364445 340509
rect 364379 340444 364380 340508
rect 364444 340444 364445 340508
rect 364379 340443 364445 340444
rect 366587 340508 366653 340509
rect 366587 340444 366588 340508
rect 366652 340444 366653 340508
rect 366587 340443 366653 340444
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 361622 266253 361682 340443
rect 361794 327454 362414 338000
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 300000 362414 326898
rect 362243 291454 362563 291486
rect 362243 291218 362285 291454
rect 362521 291218 362563 291454
rect 362243 291134 362563 291218
rect 362243 290898 362285 291134
rect 362521 290898 362563 291134
rect 362243 290866 362563 290898
rect 363541 273454 363861 273486
rect 363541 273218 363583 273454
rect 363819 273218 363861 273454
rect 363541 273134 363861 273218
rect 363541 272898 363583 273134
rect 363819 272898 363861 273134
rect 363541 272866 363861 272898
rect 361619 266252 361685 266253
rect 361619 266188 361620 266252
rect 361684 266188 361685 266252
rect 361619 266187 361685 266188
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 361622 194581 361682 266187
rect 361794 255454 362414 266000
rect 364382 265845 364442 340443
rect 368246 339510 368306 368430
rect 368246 339450 368490 339510
rect 365514 331174 366134 338000
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 300000 366134 330618
rect 368430 296730 368490 339450
rect 369234 334894 369854 338000
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 300000 369854 334338
rect 368430 296670 369410 296730
rect 364840 291454 365160 291486
rect 364840 291218 364882 291454
rect 365118 291218 365160 291454
rect 364840 291134 365160 291218
rect 364840 290898 364882 291134
rect 365118 290898 365160 291134
rect 364840 290866 365160 290898
rect 367437 291454 367757 291486
rect 367437 291218 367479 291454
rect 367715 291218 367757 291454
rect 367437 291134 367757 291218
rect 367437 290898 367479 291134
rect 367715 290898 367757 291134
rect 367437 290866 367757 290898
rect 369350 283933 369410 296670
rect 371190 295085 371250 438907
rect 371374 298077 371434 439451
rect 371558 438973 371618 582931
rect 371739 572252 371805 572253
rect 371739 572188 371740 572252
rect 371804 572188 371805 572252
rect 371739 572187 371805 572188
rect 371555 438972 371621 438973
rect 371555 438908 371556 438972
rect 371620 438908 371621 438972
rect 371555 438907 371621 438908
rect 371742 428229 371802 572187
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372475 439108 372541 439109
rect 372475 439044 372476 439108
rect 372540 439044 372541 439108
rect 372475 439043 372541 439044
rect 371923 428772 371989 428773
rect 371923 428708 371924 428772
rect 371988 428708 371989 428772
rect 371923 428707 371989 428708
rect 371739 428228 371805 428229
rect 371739 428164 371740 428228
rect 371804 428164 371805 428228
rect 371739 428163 371805 428164
rect 371371 298076 371437 298077
rect 371371 298012 371372 298076
rect 371436 298012 371437 298076
rect 371371 298011 371437 298012
rect 371742 295357 371802 428163
rect 371926 298077 371986 428707
rect 371923 298076 371989 298077
rect 371923 298012 371924 298076
rect 371988 298012 371989 298076
rect 371923 298011 371989 298012
rect 372478 296173 372538 439043
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372475 296172 372541 296173
rect 372475 296108 372476 296172
rect 372540 296108 372541 296172
rect 372475 296107 372541 296108
rect 371555 295356 371621 295357
rect 371555 295292 371556 295356
rect 371620 295292 371621 295356
rect 371555 295291 371621 295292
rect 371739 295356 371805 295357
rect 371739 295292 371740 295356
rect 371804 295292 371805 295356
rect 371739 295291 371805 295292
rect 371187 295084 371253 295085
rect 371187 295020 371188 295084
rect 371252 295020 371253 295084
rect 371187 295019 371253 295020
rect 369347 283932 369413 283933
rect 369347 283868 369348 283932
rect 369412 283868 369413 283932
rect 369347 283867 369413 283868
rect 366138 273454 366458 273486
rect 366138 273218 366180 273454
rect 366416 273218 366458 273454
rect 366138 273134 366458 273218
rect 366138 272898 366180 273134
rect 366416 272898 366458 273134
rect 366138 272866 366458 272898
rect 364379 265844 364445 265845
rect 364379 265780 364380 265844
rect 364444 265780 364445 265844
rect 364379 265779 364445 265780
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 228000 362414 254898
rect 364382 248430 364442 265779
rect 365514 259174 366134 266000
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 364382 248370 364810 248430
rect 364750 233250 364810 248370
rect 364750 233190 365178 233250
rect 365118 225725 365178 233190
rect 365514 228000 366134 258618
rect 369234 262894 369854 266000
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 228000 369854 262338
rect 365115 225724 365181 225725
rect 365115 225660 365116 225724
rect 365180 225660 365181 225724
rect 365115 225659 365181 225660
rect 366587 225724 366653 225725
rect 366587 225660 366588 225724
rect 366652 225660 366653 225724
rect 366587 225659 366653 225660
rect 362243 219454 362563 219486
rect 362243 219218 362285 219454
rect 362521 219218 362563 219454
rect 362243 219134 362563 219218
rect 362243 218898 362285 219134
rect 362521 218898 362563 219134
rect 362243 218866 362563 218898
rect 364840 219454 365160 219486
rect 364840 219218 364882 219454
rect 365118 219218 365160 219454
rect 364840 219134 365160 219218
rect 364840 218898 364882 219134
rect 365118 218898 365160 219134
rect 364840 218866 365160 218898
rect 363541 201454 363861 201486
rect 363541 201218 363583 201454
rect 363819 201218 363861 201454
rect 363541 201134 363861 201218
rect 363541 200898 363583 201134
rect 363819 200898 363861 201134
rect 363541 200866 363861 200898
rect 366138 201454 366458 201486
rect 366138 201218 366180 201454
rect 366416 201218 366458 201454
rect 366138 201134 366458 201218
rect 366138 200898 366180 201134
rect 366416 200898 366458 201134
rect 366138 200866 366458 200898
rect 366590 196485 366650 225659
rect 367437 219454 367757 219486
rect 367437 219218 367479 219454
rect 367715 219218 367757 219454
rect 367437 219134 367757 219218
rect 367437 218898 367479 219134
rect 367715 218898 367757 219134
rect 367437 218866 367757 218898
rect 365299 196484 365365 196485
rect 365299 196420 365300 196484
rect 365364 196420 365365 196484
rect 365299 196419 365365 196420
rect 366587 196484 366653 196485
rect 366587 196420 366588 196484
rect 366652 196420 366653 196484
rect 366587 196419 366653 196420
rect 361619 194580 361685 194581
rect 361619 194516 361620 194580
rect 361684 194516 361685 194580
rect 361619 194515 361685 194516
rect 362723 194580 362789 194581
rect 362723 194516 362724 194580
rect 362788 194516 362789 194580
rect 362723 194515 362789 194516
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 361794 183454 362414 194000
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 156000 362414 182898
rect 362243 147454 362563 147486
rect 362243 147218 362285 147454
rect 362521 147218 362563 147454
rect 362243 147134 362563 147218
rect 362243 146898 362285 147134
rect 362521 146898 362563 147134
rect 362243 146866 362563 146898
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 362726 123997 362786 194515
rect 364840 147454 365160 147486
rect 364840 147218 364882 147454
rect 365118 147218 365160 147454
rect 364840 147134 365160 147218
rect 364840 146898 364882 147134
rect 365118 146898 365160 147134
rect 364840 146866 365160 146898
rect 363541 129454 363861 129486
rect 363541 129218 363583 129454
rect 363819 129218 363861 129454
rect 363541 129134 363861 129218
rect 363541 128898 363583 129134
rect 363819 128898 363861 129134
rect 363541 128866 363861 128898
rect 365302 123997 365362 196419
rect 365514 187174 366134 194000
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 156000 366134 186618
rect 369234 190894 369854 194000
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 156000 369854 190338
rect 371187 152964 371253 152965
rect 371187 152900 371188 152964
rect 371252 152900 371253 152964
rect 371187 152899 371253 152900
rect 371190 148341 371250 152899
rect 371558 152693 371618 295291
rect 372478 294130 372538 296107
rect 371926 294070 372538 294130
rect 371926 277410 371986 294070
rect 372291 289916 372357 289917
rect 372291 289852 372292 289916
rect 372356 289852 372357 289916
rect 372291 289851 372357 289852
rect 372107 289508 372173 289509
rect 372107 289444 372108 289508
rect 372172 289444 372173 289508
rect 372107 289443 372173 289444
rect 371742 277350 371986 277410
rect 371555 152692 371621 152693
rect 371555 152628 371556 152692
rect 371620 152628 371621 152692
rect 371555 152627 371621 152628
rect 371742 152149 371802 277350
rect 371923 269924 371989 269925
rect 371923 269860 371924 269924
rect 371988 269860 371989 269924
rect 371923 269859 371989 269860
rect 371926 203557 371986 269859
rect 372110 231709 372170 289443
rect 372294 231845 372354 289851
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372291 231844 372357 231845
rect 372291 231780 372292 231844
rect 372356 231780 372357 231844
rect 372291 231779 372357 231780
rect 372107 231708 372173 231709
rect 372107 231644 372108 231708
rect 372172 231644 372173 231708
rect 372107 231643 372173 231644
rect 371923 203556 371989 203557
rect 371923 203492 371924 203556
rect 371988 203492 371989 203556
rect 371923 203491 371989 203492
rect 371923 158812 371989 158813
rect 371923 158748 371924 158812
rect 371988 158748 371989 158812
rect 371923 158747 371989 158748
rect 371739 152148 371805 152149
rect 371739 152084 371740 152148
rect 371804 152084 371805 152148
rect 371739 152083 371805 152084
rect 371187 148340 371253 148341
rect 371187 148276 371188 148340
rect 371252 148276 371253 148340
rect 371187 148275 371253 148276
rect 367437 147454 367757 147486
rect 367437 147218 367479 147454
rect 367715 147218 367757 147454
rect 367437 147134 367757 147218
rect 367437 146898 367479 147134
rect 367715 146898 367757 147134
rect 367437 146866 367757 146898
rect 366138 129454 366458 129486
rect 366138 129218 366180 129454
rect 366416 129218 366458 129454
rect 366138 129134 366458 129218
rect 366138 128898 366180 129134
rect 366416 128898 366458 129134
rect 366138 128866 366458 128898
rect 371926 127397 371986 158747
rect 372110 153781 372170 231643
rect 372107 153780 372173 153781
rect 372107 153716 372108 153780
rect 372172 153716 372173 153780
rect 372107 153715 372173 153716
rect 372294 153237 372354 231779
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372291 153236 372357 153237
rect 372291 153172 372292 153236
rect 372356 153172 372357 153236
rect 372291 153171 372357 153172
rect 371923 127396 371989 127397
rect 371923 127332 371924 127396
rect 371988 127332 371989 127396
rect 371923 127331 371989 127332
rect 362723 123996 362789 123997
rect 362723 123932 362724 123996
rect 362788 123932 362789 123996
rect 362723 123931 362789 123932
rect 365299 123996 365365 123997
rect 365299 123932 365300 123996
rect 365364 123932 365365 123996
rect 365299 123931 365365 123932
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 111454 362414 122000
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 115174 366134 122000
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 118894 369854 122000
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 588000 434414 614898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 588000 438134 618618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 588000 441854 622338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 434243 579454 434563 579486
rect 434243 579218 434285 579454
rect 434521 579218 434563 579454
rect 434243 579134 434563 579218
rect 434243 578898 434285 579134
rect 434521 578898 434563 579134
rect 434243 578866 434563 578898
rect 436840 579454 437160 579486
rect 436840 579218 436882 579454
rect 437118 579218 437160 579454
rect 436840 579134 437160 579218
rect 436840 578898 436882 579134
rect 437118 578898 437160 579134
rect 436840 578866 437160 578898
rect 439437 579454 439757 579486
rect 439437 579218 439479 579454
rect 439715 579218 439757 579454
rect 439437 579134 439757 579218
rect 439437 578898 439479 579134
rect 439715 578898 439757 579134
rect 439437 578866 439757 578898
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 435541 561454 435861 561486
rect 435541 561218 435583 561454
rect 435819 561218 435861 561454
rect 435541 561134 435861 561218
rect 435541 560898 435583 561134
rect 435819 560898 435861 561134
rect 435541 560866 435861 560898
rect 438138 561454 438458 561486
rect 438138 561218 438180 561454
rect 438416 561218 438458 561454
rect 438138 561134 438458 561218
rect 438138 560898 438180 561134
rect 438416 560898 438458 561134
rect 438138 560866 438458 560898
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 433794 543454 434414 554000
rect 435219 553484 435285 553485
rect 435219 553420 435220 553484
rect 435284 553420 435285 553484
rect 435219 553419 435285 553420
rect 436691 553484 436757 553485
rect 436691 553420 436692 553484
rect 436756 553420 436757 553484
rect 436691 553419 436757 553420
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 516000 434414 542898
rect 434243 507454 434563 507486
rect 434243 507218 434285 507454
rect 434521 507218 434563 507454
rect 434243 507134 434563 507218
rect 434243 506898 434285 507134
rect 434521 506898 434563 507134
rect 434243 506866 434563 506898
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 435222 483989 435282 553419
rect 435541 489454 435861 489486
rect 435541 489218 435583 489454
rect 435819 489218 435861 489454
rect 435541 489134 435861 489218
rect 435541 488898 435583 489134
rect 435819 488898 435861 489134
rect 435541 488866 435861 488898
rect 436694 483989 436754 553419
rect 437514 547174 438134 554000
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 516000 438134 546618
rect 441234 550894 441854 554000
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 516000 441854 550338
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444603 511596 444669 511597
rect 444603 511532 444604 511596
rect 444668 511532 444669 511596
rect 444603 511531 444669 511532
rect 436840 507454 437160 507486
rect 436840 507218 436882 507454
rect 437118 507218 437160 507454
rect 436840 507134 437160 507218
rect 436840 506898 436882 507134
rect 437118 506898 437160 507134
rect 436840 506866 437160 506898
rect 439437 507454 439757 507486
rect 439437 507218 439479 507454
rect 439715 507218 439757 507454
rect 439437 507134 439757 507218
rect 439437 506898 439479 507134
rect 439715 506898 439757 507134
rect 439437 506866 439757 506898
rect 444419 500308 444485 500309
rect 444419 500244 444420 500308
rect 444484 500244 444485 500308
rect 444419 500243 444485 500244
rect 438138 489454 438458 489486
rect 438138 489218 438180 489454
rect 438416 489218 438458 489454
rect 438138 489134 438458 489218
rect 438138 488898 438180 489134
rect 438416 488898 438458 489134
rect 438138 488866 438458 488898
rect 435219 483988 435285 483989
rect 435219 483924 435220 483988
rect 435284 483924 435285 483988
rect 435219 483923 435285 483924
rect 436691 483988 436757 483989
rect 436691 483924 436692 483988
rect 436756 483924 436757 483988
rect 436691 483923 436757 483924
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 433794 471454 434414 482000
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 444000 434414 470898
rect 437514 475174 438134 482000
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444000 438134 474618
rect 441234 478894 441854 482000
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 444000 441854 478338
rect 434243 435454 434563 435486
rect 434243 435218 434285 435454
rect 434521 435218 434563 435454
rect 434243 435134 434563 435218
rect 434243 434898 434285 435134
rect 434521 434898 434563 435134
rect 434243 434866 434563 434898
rect 436840 435454 437160 435486
rect 436840 435218 436882 435454
rect 437118 435218 437160 435454
rect 436840 435134 437160 435218
rect 436840 434898 436882 435134
rect 437118 434898 437160 435134
rect 436840 434866 437160 434898
rect 439437 435454 439757 435486
rect 439437 435218 439479 435454
rect 439715 435218 439757 435454
rect 439437 435134 439757 435218
rect 439437 434898 439479 435134
rect 439715 434898 439757 435134
rect 439437 434866 439757 434898
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 435541 417454 435861 417486
rect 435541 417218 435583 417454
rect 435819 417218 435861 417454
rect 435541 417134 435861 417218
rect 435541 416898 435583 417134
rect 435819 416898 435861 417134
rect 435541 416866 435861 416898
rect 438138 417454 438458 417486
rect 438138 417218 438180 417454
rect 438416 417218 438458 417454
rect 438138 417134 438458 417218
rect 438138 416898 438180 417134
rect 438416 416898 438458 417134
rect 438138 416866 438458 416898
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 433794 399454 434414 410000
rect 434851 408644 434917 408645
rect 434851 408580 434852 408644
rect 434916 408580 434917 408644
rect 434851 408579 434917 408580
rect 436139 408644 436205 408645
rect 436139 408580 436140 408644
rect 436204 408580 436205 408644
rect 436139 408579 436205 408580
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 372000 434414 398898
rect 434243 363454 434563 363486
rect 434243 363218 434285 363454
rect 434521 363218 434563 363454
rect 434243 363134 434563 363218
rect 434243 362898 434285 363134
rect 434521 362898 434563 363134
rect 434243 362866 434563 362898
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 434854 339965 434914 408579
rect 435541 345454 435861 345486
rect 435541 345218 435583 345454
rect 435819 345218 435861 345454
rect 435541 345134 435861 345218
rect 435541 344898 435583 345134
rect 435819 344898 435861 345134
rect 435541 344866 435861 344898
rect 436142 340101 436202 408579
rect 437514 403174 438134 410000
rect 440739 409596 440805 409597
rect 440739 409532 440740 409596
rect 440804 409532 440805 409596
rect 440739 409531 440805 409532
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 372000 438134 402618
rect 436840 363454 437160 363486
rect 436840 363218 436882 363454
rect 437118 363218 437160 363454
rect 436840 363134 437160 363218
rect 436840 362898 436882 363134
rect 437118 362898 437160 363134
rect 436840 362866 437160 362898
rect 439437 363454 439757 363486
rect 439437 363218 439479 363454
rect 439715 363218 439757 363454
rect 439437 363134 439757 363218
rect 439437 362898 439479 363134
rect 439715 362898 439757 363134
rect 439437 362866 439757 362898
rect 438138 345454 438458 345486
rect 438138 345218 438180 345454
rect 438416 345218 438458 345454
rect 438138 345134 438458 345218
rect 438138 344898 438180 345134
rect 438416 344898 438458 345134
rect 438138 344866 438458 344898
rect 440742 340101 440802 409531
rect 441234 406894 441854 410000
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 372000 441854 406338
rect 444422 357237 444482 500243
rect 444606 367573 444666 511531
rect 444787 500852 444853 500853
rect 444787 500788 444788 500852
rect 444852 500788 444853 500852
rect 444787 500787 444853 500788
rect 444603 367572 444669 367573
rect 444603 367508 444604 367572
rect 444668 367508 444669 367572
rect 444603 367507 444669 367508
rect 444790 364350 444850 500787
rect 444606 364290 444850 364350
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444419 357236 444485 357237
rect 444419 357172 444420 357236
rect 444484 357172 444485 357236
rect 444419 357171 444485 357172
rect 444422 356285 444482 357171
rect 444606 356829 444666 364290
rect 444603 356828 444669 356829
rect 444603 356764 444604 356828
rect 444668 356764 444669 356828
rect 444603 356763 444669 356764
rect 444419 356284 444485 356285
rect 444419 356220 444420 356284
rect 444484 356220 444485 356284
rect 444419 356219 444485 356220
rect 436139 340100 436205 340101
rect 436139 340036 436140 340100
rect 436204 340036 436205 340100
rect 436139 340035 436205 340036
rect 440739 340100 440805 340101
rect 440739 340036 440740 340100
rect 440804 340036 440805 340100
rect 440739 340035 440805 340036
rect 434851 339964 434917 339965
rect 434851 339900 434852 339964
rect 434916 339900 434917 339964
rect 434851 339899 434917 339900
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 433794 327454 434414 338000
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 300000 434414 326898
rect 437514 331174 438134 338000
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 300000 438134 330618
rect 441234 334894 441854 338000
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 300000 441854 334338
rect 434243 291454 434563 291486
rect 434243 291218 434285 291454
rect 434521 291218 434563 291454
rect 434243 291134 434563 291218
rect 434243 290898 434285 291134
rect 434521 290898 434563 291134
rect 434243 290866 434563 290898
rect 436840 291454 437160 291486
rect 436840 291218 436882 291454
rect 437118 291218 437160 291454
rect 436840 291134 437160 291218
rect 436840 290898 436882 291134
rect 437118 290898 437160 291134
rect 436840 290866 437160 290898
rect 439437 291454 439757 291486
rect 439437 291218 439479 291454
rect 439715 291218 439757 291454
rect 439437 291134 439757 291218
rect 439437 290898 439479 291134
rect 439715 290898 439757 291134
rect 439437 290866 439757 290898
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 435541 273454 435861 273486
rect 435541 273218 435583 273454
rect 435819 273218 435861 273454
rect 435541 273134 435861 273218
rect 435541 272898 435583 273134
rect 435819 272898 435861 273134
rect 435541 272866 435861 272898
rect 438138 273454 438458 273486
rect 438138 273218 438180 273454
rect 438416 273218 438458 273454
rect 438138 273134 438458 273218
rect 438138 272898 438180 273134
rect 438416 272898 438458 273134
rect 438138 272866 438458 272898
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 433794 255454 434414 266000
rect 436691 265572 436757 265573
rect 436691 265508 436692 265572
rect 436756 265508 436757 265572
rect 436691 265507 436757 265508
rect 435219 265028 435285 265029
rect 435219 264964 435220 265028
rect 435284 264964 435285 265028
rect 435219 264963 435285 264964
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 228000 434414 254898
rect 434243 219454 434563 219486
rect 434243 219218 434285 219454
rect 434521 219218 434563 219454
rect 434243 219134 434563 219218
rect 434243 218898 434285 219134
rect 434521 218898 434563 219134
rect 434243 218866 434563 218898
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 435222 196077 435282 264963
rect 435541 201454 435861 201486
rect 435541 201218 435583 201454
rect 435819 201218 435861 201454
rect 435541 201134 435861 201218
rect 435541 200898 435583 201134
rect 435819 200898 435861 201134
rect 435541 200866 435861 200898
rect 436694 196077 436754 265507
rect 437514 259174 438134 266000
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 228000 438134 258618
rect 441234 262894 441854 266000
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 228000 441854 262338
rect 436840 219454 437160 219486
rect 436840 219218 436882 219454
rect 437118 219218 437160 219454
rect 436840 219134 437160 219218
rect 436840 218898 436882 219134
rect 437118 218898 437160 219134
rect 436840 218866 437160 218898
rect 439437 219454 439757 219486
rect 439437 219218 439479 219454
rect 439715 219218 439757 219454
rect 439437 219134 439757 219218
rect 439437 218898 439479 219134
rect 439715 218898 439757 219134
rect 439437 218866 439757 218898
rect 444422 212261 444482 356219
rect 444606 267749 444666 356763
rect 444787 354652 444853 354653
rect 444787 354588 444788 354652
rect 444852 354588 444853 354652
rect 444787 354587 444853 354588
rect 444603 267748 444669 267749
rect 444603 267684 444604 267748
rect 444668 267684 444669 267748
rect 444603 267683 444669 267684
rect 444606 212805 444666 267683
rect 444603 212804 444669 212805
rect 444603 212740 444604 212804
rect 444668 212740 444669 212804
rect 444603 212739 444669 212740
rect 444790 212397 444850 354587
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444787 212396 444853 212397
rect 444787 212332 444788 212396
rect 444852 212332 444853 212396
rect 444787 212331 444853 212332
rect 444419 212260 444485 212261
rect 444419 212196 444420 212260
rect 444484 212196 444485 212260
rect 444419 212195 444485 212196
rect 444790 211173 444850 212331
rect 444787 211172 444853 211173
rect 444787 211108 444788 211172
rect 444852 211108 444853 211172
rect 444787 211107 444853 211108
rect 438138 201454 438458 201486
rect 438138 201218 438180 201454
rect 438416 201218 438458 201454
rect 438138 201134 438458 201218
rect 444419 201244 444485 201245
rect 444419 201180 444420 201244
rect 444484 201180 444485 201244
rect 444419 201179 444485 201180
rect 438138 200898 438180 201134
rect 438416 200898 438458 201134
rect 438138 200866 438458 200898
rect 435219 196076 435285 196077
rect 435219 196012 435220 196076
rect 435284 196012 435285 196076
rect 435219 196011 435285 196012
rect 436691 196076 436757 196077
rect 436691 196012 436692 196076
rect 436756 196012 436757 196076
rect 436691 196011 436757 196012
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 433794 183454 434414 194000
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 156000 434414 182898
rect 437514 187174 438134 194000
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 156000 438134 186618
rect 441234 190894 441854 194000
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 156000 441854 190338
rect 434243 147454 434563 147486
rect 434243 147218 434285 147454
rect 434521 147218 434563 147454
rect 434243 147134 434563 147218
rect 434243 146898 434285 147134
rect 434521 146898 434563 147134
rect 434243 146866 434563 146898
rect 436840 147454 437160 147486
rect 436840 147218 436882 147454
rect 437118 147218 437160 147454
rect 436840 147134 437160 147218
rect 436840 146898 436882 147134
rect 437118 146898 437160 147134
rect 436840 146866 437160 146898
rect 439437 147454 439757 147486
rect 439437 147218 439479 147454
rect 439715 147218 439757 147454
rect 439437 147134 439757 147218
rect 439437 146898 439479 147134
rect 439715 146898 439757 147134
rect 439437 146866 439757 146898
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 444422 135013 444482 201179
rect 444603 198932 444669 198933
rect 444603 198868 444604 198932
rect 444668 198868 444669 198932
rect 444603 198867 444669 198868
rect 444606 158813 444666 198867
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444787 169692 444853 169693
rect 444787 169628 444788 169692
rect 444852 169628 444853 169692
rect 444787 169627 444853 169628
rect 444790 169013 444850 169627
rect 444787 169012 444853 169013
rect 444787 168948 444788 169012
rect 444852 168948 444853 169012
rect 444787 168947 444853 168948
rect 444603 158812 444669 158813
rect 444603 158748 444604 158812
rect 444668 158748 444669 158812
rect 444603 158747 444669 158748
rect 444790 156501 444850 168947
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444787 156500 444853 156501
rect 444787 156436 444788 156500
rect 444852 156436 444853 156500
rect 444787 156435 444853 156436
rect 444419 135012 444485 135013
rect 444419 134948 444420 135012
rect 444484 134948 444485 135012
rect 444419 134947 444485 134948
rect 435541 129454 435861 129486
rect 435541 129218 435583 129454
rect 435819 129218 435861 129454
rect 435541 129134 435861 129218
rect 435541 128898 435583 129134
rect 435819 128898 435861 129134
rect 435541 128866 435861 128898
rect 438138 129454 438458 129486
rect 438138 129218 438180 129454
rect 438416 129218 438458 129454
rect 438138 129134 438458 129218
rect 438138 128898 438180 129134
rect 438416 128898 438458 129134
rect 438138 128866 438458 128898
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 111454 434414 122000
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 115174 438134 122000
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 118894 441854 122000
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 588000 506414 614898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 588000 510134 618618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 588000 513854 622338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 506243 579454 506563 579486
rect 506243 579218 506285 579454
rect 506521 579218 506563 579454
rect 506243 579134 506563 579218
rect 506243 578898 506285 579134
rect 506521 578898 506563 579134
rect 506243 578866 506563 578898
rect 508840 579454 509160 579486
rect 508840 579218 508882 579454
rect 509118 579218 509160 579454
rect 508840 579134 509160 579218
rect 508840 578898 508882 579134
rect 509118 578898 509160 579134
rect 508840 578866 509160 578898
rect 511437 579454 511757 579486
rect 511437 579218 511479 579454
rect 511715 579218 511757 579454
rect 511437 579134 511757 579218
rect 511437 578898 511479 579134
rect 511715 578898 511757 579134
rect 511437 578866 511757 578898
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 507541 561454 507861 561486
rect 507541 561218 507583 561454
rect 507819 561218 507861 561454
rect 507541 561134 507861 561218
rect 507541 560898 507583 561134
rect 507819 560898 507861 561134
rect 507541 560866 507861 560898
rect 510138 561454 510458 561486
rect 510138 561218 510180 561454
rect 510416 561218 510458 561454
rect 510138 561134 510458 561218
rect 510138 560898 510180 561134
rect 510416 560898 510458 561134
rect 510138 560866 510458 560898
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 505794 543454 506414 554000
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 516000 506414 542898
rect 509514 547174 510134 554000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 516000 510134 546618
rect 513234 550894 513854 554000
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 516000 513854 550338
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 506243 507454 506563 507486
rect 506243 507218 506285 507454
rect 506521 507218 506563 507454
rect 506243 507134 506563 507218
rect 506243 506898 506285 507134
rect 506521 506898 506563 507134
rect 506243 506866 506563 506898
rect 508840 507454 509160 507486
rect 508840 507218 508882 507454
rect 509118 507218 509160 507454
rect 508840 507134 509160 507218
rect 508840 506898 508882 507134
rect 509118 506898 509160 507134
rect 508840 506866 509160 506898
rect 511437 507454 511757 507486
rect 511437 507218 511479 507454
rect 511715 507218 511757 507454
rect 511437 507134 511757 507218
rect 511437 506898 511479 507134
rect 511715 506898 511757 507134
rect 511437 506866 511757 506898
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 507541 489454 507861 489486
rect 507541 489218 507583 489454
rect 507819 489218 507861 489454
rect 507541 489134 507861 489218
rect 507541 488898 507583 489134
rect 507819 488898 507861 489134
rect 507541 488866 507861 488898
rect 510138 489454 510458 489486
rect 510138 489218 510180 489454
rect 510416 489218 510458 489454
rect 510138 489134 510458 489218
rect 510138 488898 510180 489134
rect 510416 488898 510458 489134
rect 510138 488866 510458 488898
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 505794 471454 506414 482000
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 444000 506414 470898
rect 509514 475174 510134 482000
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 444000 510134 474618
rect 513234 478894 513854 482000
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 444000 513854 478338
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516179 439516 516245 439517
rect 516179 439452 516180 439516
rect 516244 439452 516245 439516
rect 516179 439451 516245 439452
rect 506243 435454 506563 435486
rect 506243 435218 506285 435454
rect 506521 435218 506563 435454
rect 506243 435134 506563 435218
rect 506243 434898 506285 435134
rect 506521 434898 506563 435134
rect 506243 434866 506563 434898
rect 508840 435454 509160 435486
rect 508840 435218 508882 435454
rect 509118 435218 509160 435454
rect 508840 435134 509160 435218
rect 508840 434898 508882 435134
rect 509118 434898 509160 435134
rect 508840 434866 509160 434898
rect 511437 435454 511757 435486
rect 511437 435218 511479 435454
rect 511715 435218 511757 435454
rect 511437 435134 511757 435218
rect 511437 434898 511479 435134
rect 511715 434898 511757 435134
rect 511437 434866 511757 434898
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 507541 417454 507861 417486
rect 507541 417218 507583 417454
rect 507819 417218 507861 417454
rect 507541 417134 507861 417218
rect 507541 416898 507583 417134
rect 507819 416898 507861 417134
rect 507541 416866 507861 416898
rect 510138 417454 510458 417486
rect 510138 417218 510180 417454
rect 510416 417218 510458 417454
rect 510138 417134 510458 417218
rect 510138 416898 510180 417134
rect 510416 416898 510458 417134
rect 510138 416866 510458 416898
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 505794 399454 506414 410000
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 372000 506414 398898
rect 509514 403174 510134 410000
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 372000 510134 402618
rect 513234 406894 513854 410000
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 372000 513854 406338
rect 506243 363454 506563 363486
rect 506243 363218 506285 363454
rect 506521 363218 506563 363454
rect 506243 363134 506563 363218
rect 506243 362898 506285 363134
rect 506521 362898 506563 363134
rect 506243 362866 506563 362898
rect 508840 363454 509160 363486
rect 508840 363218 508882 363454
rect 509118 363218 509160 363454
rect 508840 363134 509160 363218
rect 508840 362898 508882 363134
rect 509118 362898 509160 363134
rect 508840 362866 509160 362898
rect 511437 363454 511757 363486
rect 511437 363218 511479 363454
rect 511715 363218 511757 363454
rect 511437 363134 511757 363218
rect 511437 362898 511479 363134
rect 511715 362898 511757 363134
rect 511437 362866 511757 362898
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 507541 345454 507861 345486
rect 507541 345218 507583 345454
rect 507819 345218 507861 345454
rect 507541 345134 507861 345218
rect 507541 344898 507583 345134
rect 507819 344898 507861 345134
rect 507541 344866 507861 344898
rect 510138 345454 510458 345486
rect 510138 345218 510180 345454
rect 510416 345218 510458 345454
rect 510138 345134 510458 345218
rect 510138 344898 510180 345134
rect 510416 344898 510458 345134
rect 510138 344866 510458 344898
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 505794 327454 506414 338000
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 300000 506414 326898
rect 509514 331174 510134 338000
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 300000 510134 330618
rect 513234 334894 513854 338000
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 300000 513854 334338
rect 516182 295901 516242 439451
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516363 298212 516429 298213
rect 516363 298148 516364 298212
rect 516428 298148 516429 298212
rect 516363 298147 516429 298148
rect 516179 295900 516245 295901
rect 516179 295836 516180 295900
rect 516244 295836 516245 295900
rect 516179 295835 516245 295836
rect 516366 293861 516426 298147
rect 516363 293860 516429 293861
rect 516363 293796 516364 293860
rect 516428 293796 516429 293860
rect 516363 293795 516429 293796
rect 506243 291454 506563 291486
rect 506243 291218 506285 291454
rect 506521 291218 506563 291454
rect 506243 291134 506563 291218
rect 506243 290898 506285 291134
rect 506521 290898 506563 291134
rect 506243 290866 506563 290898
rect 508840 291454 509160 291486
rect 508840 291218 508882 291454
rect 509118 291218 509160 291454
rect 508840 291134 509160 291218
rect 508840 290898 508882 291134
rect 509118 290898 509160 291134
rect 508840 290866 509160 290898
rect 511437 291454 511757 291486
rect 511437 291218 511479 291454
rect 511715 291218 511757 291454
rect 511437 291134 511757 291218
rect 511437 290898 511479 291134
rect 511715 290898 511757 291134
rect 511437 290866 511757 290898
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 507541 273454 507861 273486
rect 507541 273218 507583 273454
rect 507819 273218 507861 273454
rect 507541 273134 507861 273218
rect 507541 272898 507583 273134
rect 507819 272898 507861 273134
rect 507541 272866 507861 272898
rect 510138 273454 510458 273486
rect 510138 273218 510180 273454
rect 510416 273218 510458 273454
rect 510138 273134 510458 273218
rect 510138 272898 510180 273134
rect 510416 272898 510458 273134
rect 510138 272866 510458 272898
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 505794 255454 506414 266000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 228000 506414 254898
rect 509514 259174 510134 266000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 228000 510134 258618
rect 513234 262894 513854 266000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 228000 513854 262338
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 506243 219454 506563 219486
rect 506243 219218 506285 219454
rect 506521 219218 506563 219454
rect 506243 219134 506563 219218
rect 506243 218898 506285 219134
rect 506521 218898 506563 219134
rect 506243 218866 506563 218898
rect 508840 219454 509160 219486
rect 508840 219218 508882 219454
rect 509118 219218 509160 219454
rect 508840 219134 509160 219218
rect 508840 218898 508882 219134
rect 509118 218898 509160 219134
rect 508840 218866 509160 218898
rect 511437 219454 511757 219486
rect 511437 219218 511479 219454
rect 511715 219218 511757 219454
rect 511437 219134 511757 219218
rect 511437 218898 511479 219134
rect 511715 218898 511757 219134
rect 511437 218866 511757 218898
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 507541 201454 507861 201486
rect 507541 201218 507583 201454
rect 507819 201218 507861 201454
rect 507541 201134 507861 201218
rect 507541 200898 507583 201134
rect 507819 200898 507861 201134
rect 507541 200866 507861 200898
rect 510138 201454 510458 201486
rect 510138 201218 510180 201454
rect 510416 201218 510458 201454
rect 510138 201134 510458 201218
rect 510138 200898 510180 201134
rect 510416 200898 510458 201134
rect 510138 200866 510458 200898
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 505794 183454 506414 194000
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 156000 506414 182898
rect 509514 187174 510134 194000
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 156000 510134 186618
rect 513234 190894 513854 194000
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 156000 513854 190338
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 514155 152964 514221 152965
rect 514155 152900 514156 152964
rect 514220 152900 514221 152964
rect 514155 152899 514221 152900
rect 513971 152420 514037 152421
rect 513971 152356 513972 152420
rect 514036 152356 514037 152420
rect 513971 152355 514037 152356
rect 513974 151333 514034 152355
rect 514158 151877 514218 152899
rect 514339 152012 514405 152013
rect 514339 151948 514340 152012
rect 514404 151948 514405 152012
rect 514339 151947 514405 151948
rect 514155 151876 514221 151877
rect 514155 151812 514156 151876
rect 514220 151812 514221 151876
rect 514155 151811 514221 151812
rect 514342 151469 514402 151947
rect 514339 151468 514405 151469
rect 514339 151404 514340 151468
rect 514404 151404 514405 151468
rect 514339 151403 514405 151404
rect 513971 151332 514037 151333
rect 513971 151268 513972 151332
rect 514036 151268 514037 151332
rect 513971 151267 514037 151268
rect 506243 147454 506563 147486
rect 506243 147218 506285 147454
rect 506521 147218 506563 147454
rect 506243 147134 506563 147218
rect 506243 146898 506285 147134
rect 506521 146898 506563 147134
rect 506243 146866 506563 146898
rect 508840 147454 509160 147486
rect 508840 147218 508882 147454
rect 509118 147218 509160 147454
rect 508840 147134 509160 147218
rect 508840 146898 508882 147134
rect 509118 146898 509160 147134
rect 508840 146866 509160 146898
rect 511437 147454 511757 147486
rect 511437 147218 511479 147454
rect 511715 147218 511757 147454
rect 511437 147134 511757 147218
rect 511437 146898 511479 147134
rect 511715 146898 511757 147134
rect 511437 146866 511757 146898
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 507541 129454 507861 129486
rect 507541 129218 507583 129454
rect 507819 129218 507861 129454
rect 507541 129134 507861 129218
rect 507541 128898 507583 129134
rect 507819 128898 507861 129134
rect 507541 128866 507861 128898
rect 510138 129454 510458 129486
rect 510138 129218 510180 129454
rect 510416 129218 510458 129454
rect 510138 129134 510458 129218
rect 510138 128898 510180 129134
rect 510416 128898 510458 129134
rect 510138 128866 510458 128898
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 111454 506414 122000
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 115174 510134 122000
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 118894 513854 122000
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 162285 183218 162521 183454
rect 162285 182898 162521 183134
rect 164882 183218 165118 183454
rect 164882 182898 165118 183134
rect 167479 183218 167715 183454
rect 167479 182898 167715 183134
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 163583 165218 163819 165454
rect 163583 164898 163819 165134
rect 166180 165218 166416 165454
rect 166180 164898 166416 165134
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 162285 147218 162521 147454
rect 162285 146898 162521 147134
rect 164882 147218 165118 147454
rect 164882 146898 165118 147134
rect 167479 147218 167715 147454
rect 167479 146898 167715 147134
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 163583 129218 163819 129454
rect 163583 128898 163819 129134
rect 166180 129218 166416 129454
rect 166180 128898 166416 129134
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 204250 291218 204486 291454
rect 204250 290898 204486 291134
rect 234970 291218 235206 291454
rect 234970 290898 235206 291134
rect 265690 291218 265926 291454
rect 265690 290898 265926 291134
rect 296410 291218 296646 291454
rect 296410 290898 296646 291134
rect 219610 273218 219846 273454
rect 219610 272898 219846 273134
rect 250330 273218 250566 273454
rect 250330 272898 250566 273134
rect 281050 273218 281286 273454
rect 281050 272898 281286 273134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 204250 255218 204486 255454
rect 204250 254898 204486 255134
rect 234970 255218 235206 255454
rect 234970 254898 235206 255134
rect 265690 255218 265926 255454
rect 265690 254898 265926 255134
rect 296410 255218 296646 255454
rect 296410 254898 296646 255134
rect 219610 237218 219846 237454
rect 219610 236898 219846 237134
rect 250330 237218 250566 237454
rect 250330 236898 250566 237134
rect 281050 237218 281286 237454
rect 281050 236898 281286 237134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 204250 219218 204486 219454
rect 204250 218898 204486 219134
rect 234970 219218 235206 219454
rect 234970 218898 235206 219134
rect 265690 219218 265926 219454
rect 265690 218898 265926 219134
rect 296410 219218 296646 219454
rect 296410 218898 296646 219134
rect 219610 201218 219846 201454
rect 219610 200898 219846 201134
rect 250330 201218 250566 201454
rect 250330 200898 250566 201134
rect 281050 201218 281286 201454
rect 281050 200898 281286 201134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 204250 183218 204486 183454
rect 204250 182898 204486 183134
rect 234970 183218 235206 183454
rect 234970 182898 235206 183134
rect 265690 183218 265926 183454
rect 265690 182898 265926 183134
rect 296410 183218 296646 183454
rect 296410 182898 296646 183134
rect 219610 165218 219846 165454
rect 219610 164898 219846 165134
rect 250330 165218 250566 165454
rect 250330 164898 250566 165134
rect 281050 165218 281286 165454
rect 281050 164898 281286 165134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 204250 147218 204486 147454
rect 204250 146898 204486 147134
rect 234970 147218 235206 147454
rect 234970 146898 235206 147134
rect 265690 147218 265926 147454
rect 265690 146898 265926 147134
rect 296410 147218 296646 147454
rect 296410 146898 296646 147134
rect 219610 129218 219846 129454
rect 219610 128898 219846 129134
rect 250330 129218 250566 129454
rect 250330 128898 250566 129134
rect 281050 129218 281286 129454
rect 281050 128898 281286 129134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 204250 111218 204486 111454
rect 204250 110898 204486 111134
rect 234970 111218 235206 111454
rect 234970 110898 235206 111134
rect 265690 111218 265926 111454
rect 265690 110898 265926 111134
rect 296410 111218 296646 111454
rect 296410 110898 296646 111134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 362285 579218 362521 579454
rect 362285 578898 362521 579134
rect 364882 579218 365118 579454
rect 364882 578898 365118 579134
rect 367479 579218 367715 579454
rect 367479 578898 367715 579134
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 363583 561218 363819 561454
rect 363583 560898 363819 561134
rect 366180 561218 366416 561454
rect 366180 560898 366416 561134
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 362285 507218 362521 507454
rect 362285 506898 362521 507134
rect 364882 507218 365118 507454
rect 364882 506898 365118 507134
rect 363583 489218 363819 489454
rect 363583 488898 363819 489134
rect 366180 489218 366416 489454
rect 366180 488898 366416 489134
rect 367479 507218 367715 507454
rect 367479 506898 367715 507134
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 362285 435218 362521 435454
rect 362285 434898 362521 435134
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 364882 435218 365118 435454
rect 364882 434898 365118 435134
rect 363583 417218 363819 417454
rect 363583 416898 363819 417134
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 367479 435218 367715 435454
rect 367479 434898 367715 435134
rect 366180 417218 366416 417454
rect 366180 416898 366416 417134
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 362285 363218 362521 363454
rect 362285 362898 362521 363134
rect 364882 363218 365118 363454
rect 364882 362898 365118 363134
rect 363583 345218 363819 345454
rect 363583 344898 363819 345134
rect 366180 345218 366416 345454
rect 366180 344898 366416 345134
rect 367479 363218 367715 363454
rect 367479 362898 367715 363134
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 362285 291218 362521 291454
rect 362285 290898 362521 291134
rect 363583 273218 363819 273454
rect 363583 272898 363819 273134
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 364882 291218 365118 291454
rect 364882 290898 365118 291134
rect 367479 291218 367715 291454
rect 367479 290898 367715 291134
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 366180 273218 366416 273454
rect 366180 272898 366416 273134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 362285 219218 362521 219454
rect 362285 218898 362521 219134
rect 364882 219218 365118 219454
rect 364882 218898 365118 219134
rect 363583 201218 363819 201454
rect 363583 200898 363819 201134
rect 366180 201218 366416 201454
rect 366180 200898 366416 201134
rect 367479 219218 367715 219454
rect 367479 218898 367715 219134
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 362285 147218 362521 147454
rect 362285 146898 362521 147134
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 364882 147218 365118 147454
rect 364882 146898 365118 147134
rect 363583 129218 363819 129454
rect 363583 128898 363819 129134
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 367479 147218 367715 147454
rect 367479 146898 367715 147134
rect 366180 129218 366416 129454
rect 366180 128898 366416 129134
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 434285 579218 434521 579454
rect 434285 578898 434521 579134
rect 436882 579218 437118 579454
rect 436882 578898 437118 579134
rect 439479 579218 439715 579454
rect 439479 578898 439715 579134
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 435583 561218 435819 561454
rect 435583 560898 435819 561134
rect 438180 561218 438416 561454
rect 438180 560898 438416 561134
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 434285 507218 434521 507454
rect 434285 506898 434521 507134
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 435583 489218 435819 489454
rect 435583 488898 435819 489134
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 436882 507218 437118 507454
rect 436882 506898 437118 507134
rect 439479 507218 439715 507454
rect 439479 506898 439715 507134
rect 438180 489218 438416 489454
rect 438180 488898 438416 489134
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 434285 435218 434521 435454
rect 434285 434898 434521 435134
rect 436882 435218 437118 435454
rect 436882 434898 437118 435134
rect 439479 435218 439715 435454
rect 439479 434898 439715 435134
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 435583 417218 435819 417454
rect 435583 416898 435819 417134
rect 438180 417218 438416 417454
rect 438180 416898 438416 417134
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 434285 363218 434521 363454
rect 434285 362898 434521 363134
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 435583 345218 435819 345454
rect 435583 344898 435819 345134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 436882 363218 437118 363454
rect 436882 362898 437118 363134
rect 439479 363218 439715 363454
rect 439479 362898 439715 363134
rect 438180 345218 438416 345454
rect 438180 344898 438416 345134
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 434285 291218 434521 291454
rect 434285 290898 434521 291134
rect 436882 291218 437118 291454
rect 436882 290898 437118 291134
rect 439479 291218 439715 291454
rect 439479 290898 439715 291134
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 435583 273218 435819 273454
rect 435583 272898 435819 273134
rect 438180 273218 438416 273454
rect 438180 272898 438416 273134
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 434285 219218 434521 219454
rect 434285 218898 434521 219134
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 435583 201218 435819 201454
rect 435583 200898 435819 201134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 436882 219218 437118 219454
rect 436882 218898 437118 219134
rect 439479 219218 439715 219454
rect 439479 218898 439715 219134
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 438180 201218 438416 201454
rect 438180 200898 438416 201134
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 434285 147218 434521 147454
rect 434285 146898 434521 147134
rect 436882 147218 437118 147454
rect 436882 146898 437118 147134
rect 439479 147218 439715 147454
rect 439479 146898 439715 147134
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 435583 129218 435819 129454
rect 435583 128898 435819 129134
rect 438180 129218 438416 129454
rect 438180 128898 438416 129134
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 506285 579218 506521 579454
rect 506285 578898 506521 579134
rect 508882 579218 509118 579454
rect 508882 578898 509118 579134
rect 511479 579218 511715 579454
rect 511479 578898 511715 579134
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 507583 561218 507819 561454
rect 507583 560898 507819 561134
rect 510180 561218 510416 561454
rect 510180 560898 510416 561134
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 506285 507218 506521 507454
rect 506285 506898 506521 507134
rect 508882 507218 509118 507454
rect 508882 506898 509118 507134
rect 511479 507218 511715 507454
rect 511479 506898 511715 507134
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 507583 489218 507819 489454
rect 507583 488898 507819 489134
rect 510180 489218 510416 489454
rect 510180 488898 510416 489134
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 506285 435218 506521 435454
rect 506285 434898 506521 435134
rect 508882 435218 509118 435454
rect 508882 434898 509118 435134
rect 511479 435218 511715 435454
rect 511479 434898 511715 435134
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 507583 417218 507819 417454
rect 507583 416898 507819 417134
rect 510180 417218 510416 417454
rect 510180 416898 510416 417134
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 506285 363218 506521 363454
rect 506285 362898 506521 363134
rect 508882 363218 509118 363454
rect 508882 362898 509118 363134
rect 511479 363218 511715 363454
rect 511479 362898 511715 363134
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 507583 345218 507819 345454
rect 507583 344898 507819 345134
rect 510180 345218 510416 345454
rect 510180 344898 510416 345134
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 506285 291218 506521 291454
rect 506285 290898 506521 291134
rect 508882 291218 509118 291454
rect 508882 290898 509118 291134
rect 511479 291218 511715 291454
rect 511479 290898 511715 291134
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 507583 273218 507819 273454
rect 507583 272898 507819 273134
rect 510180 273218 510416 273454
rect 510180 272898 510416 273134
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 506285 219218 506521 219454
rect 506285 218898 506521 219134
rect 508882 219218 509118 219454
rect 508882 218898 509118 219134
rect 511479 219218 511715 219454
rect 511479 218898 511715 219134
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 507583 201218 507819 201454
rect 507583 200898 507819 201134
rect 510180 201218 510416 201454
rect 510180 200898 510416 201134
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 506285 147218 506521 147454
rect 506285 146898 506521 147134
rect 508882 147218 509118 147454
rect 508882 146898 509118 147134
rect 511479 147218 511715 147454
rect 511479 146898 511715 147134
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 507583 129218 507819 129454
rect 507583 128898 507819 129134
rect 510180 129218 510416 129454
rect 510180 128898 510416 129134
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 362285 579454
rect 362521 579218 364882 579454
rect 365118 579218 367479 579454
rect 367715 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 434285 579454
rect 434521 579218 436882 579454
rect 437118 579218 439479 579454
rect 439715 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 506285 579454
rect 506521 579218 508882 579454
rect 509118 579218 511479 579454
rect 511715 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 362285 579134
rect 362521 578898 364882 579134
rect 365118 578898 367479 579134
rect 367715 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 434285 579134
rect 434521 578898 436882 579134
rect 437118 578898 439479 579134
rect 439715 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 506285 579134
rect 506521 578898 508882 579134
rect 509118 578898 511479 579134
rect 511715 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 363583 561454
rect 363819 561218 366180 561454
rect 366416 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 435583 561454
rect 435819 561218 438180 561454
rect 438416 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 507583 561454
rect 507819 561218 510180 561454
rect 510416 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 363583 561134
rect 363819 560898 366180 561134
rect 366416 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 435583 561134
rect 435819 560898 438180 561134
rect 438416 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 507583 561134
rect 507819 560898 510180 561134
rect 510416 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 362285 507454
rect 362521 507218 364882 507454
rect 365118 507218 367479 507454
rect 367715 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 434285 507454
rect 434521 507218 436882 507454
rect 437118 507218 439479 507454
rect 439715 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 506285 507454
rect 506521 507218 508882 507454
rect 509118 507218 511479 507454
rect 511715 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 362285 507134
rect 362521 506898 364882 507134
rect 365118 506898 367479 507134
rect 367715 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 434285 507134
rect 434521 506898 436882 507134
rect 437118 506898 439479 507134
rect 439715 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 506285 507134
rect 506521 506898 508882 507134
rect 509118 506898 511479 507134
rect 511715 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 363583 489454
rect 363819 489218 366180 489454
rect 366416 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 435583 489454
rect 435819 489218 438180 489454
rect 438416 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 507583 489454
rect 507819 489218 510180 489454
rect 510416 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 363583 489134
rect 363819 488898 366180 489134
rect 366416 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 435583 489134
rect 435819 488898 438180 489134
rect 438416 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 507583 489134
rect 507819 488898 510180 489134
rect 510416 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 362285 435454
rect 362521 435218 364882 435454
rect 365118 435218 367479 435454
rect 367715 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 434285 435454
rect 434521 435218 436882 435454
rect 437118 435218 439479 435454
rect 439715 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 506285 435454
rect 506521 435218 508882 435454
rect 509118 435218 511479 435454
rect 511715 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 362285 435134
rect 362521 434898 364882 435134
rect 365118 434898 367479 435134
rect 367715 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 434285 435134
rect 434521 434898 436882 435134
rect 437118 434898 439479 435134
rect 439715 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 506285 435134
rect 506521 434898 508882 435134
rect 509118 434898 511479 435134
rect 511715 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 363583 417454
rect 363819 417218 366180 417454
rect 366416 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 435583 417454
rect 435819 417218 438180 417454
rect 438416 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 507583 417454
rect 507819 417218 510180 417454
rect 510416 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 363583 417134
rect 363819 416898 366180 417134
rect 366416 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 435583 417134
rect 435819 416898 438180 417134
rect 438416 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 507583 417134
rect 507819 416898 510180 417134
rect 510416 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 362285 363454
rect 362521 363218 364882 363454
rect 365118 363218 367479 363454
rect 367715 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 434285 363454
rect 434521 363218 436882 363454
rect 437118 363218 439479 363454
rect 439715 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 506285 363454
rect 506521 363218 508882 363454
rect 509118 363218 511479 363454
rect 511715 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 362285 363134
rect 362521 362898 364882 363134
rect 365118 362898 367479 363134
rect 367715 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 434285 363134
rect 434521 362898 436882 363134
rect 437118 362898 439479 363134
rect 439715 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 506285 363134
rect 506521 362898 508882 363134
rect 509118 362898 511479 363134
rect 511715 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 363583 345454
rect 363819 345218 366180 345454
rect 366416 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 435583 345454
rect 435819 345218 438180 345454
rect 438416 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 507583 345454
rect 507819 345218 510180 345454
rect 510416 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 363583 345134
rect 363819 344898 366180 345134
rect 366416 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 435583 345134
rect 435819 344898 438180 345134
rect 438416 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 507583 345134
rect 507819 344898 510180 345134
rect 510416 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 204250 291454
rect 204486 291218 234970 291454
rect 235206 291218 265690 291454
rect 265926 291218 296410 291454
rect 296646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 362285 291454
rect 362521 291218 364882 291454
rect 365118 291218 367479 291454
rect 367715 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 434285 291454
rect 434521 291218 436882 291454
rect 437118 291218 439479 291454
rect 439715 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 506285 291454
rect 506521 291218 508882 291454
rect 509118 291218 511479 291454
rect 511715 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 204250 291134
rect 204486 290898 234970 291134
rect 235206 290898 265690 291134
rect 265926 290898 296410 291134
rect 296646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 362285 291134
rect 362521 290898 364882 291134
rect 365118 290898 367479 291134
rect 367715 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 434285 291134
rect 434521 290898 436882 291134
rect 437118 290898 439479 291134
rect 439715 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 506285 291134
rect 506521 290898 508882 291134
rect 509118 290898 511479 291134
rect 511715 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219610 273454
rect 219846 273218 250330 273454
rect 250566 273218 281050 273454
rect 281286 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 363583 273454
rect 363819 273218 366180 273454
rect 366416 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 435583 273454
rect 435819 273218 438180 273454
rect 438416 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 507583 273454
rect 507819 273218 510180 273454
rect 510416 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219610 273134
rect 219846 272898 250330 273134
rect 250566 272898 281050 273134
rect 281286 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 363583 273134
rect 363819 272898 366180 273134
rect 366416 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 435583 273134
rect 435819 272898 438180 273134
rect 438416 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 507583 273134
rect 507819 272898 510180 273134
rect 510416 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204250 255454
rect 204486 255218 234970 255454
rect 235206 255218 265690 255454
rect 265926 255218 296410 255454
rect 296646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204250 255134
rect 204486 254898 234970 255134
rect 235206 254898 265690 255134
rect 265926 254898 296410 255134
rect 296646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 219610 237454
rect 219846 237218 250330 237454
rect 250566 237218 281050 237454
rect 281286 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 219610 237134
rect 219846 236898 250330 237134
rect 250566 236898 281050 237134
rect 281286 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 204250 219454
rect 204486 219218 234970 219454
rect 235206 219218 265690 219454
rect 265926 219218 296410 219454
rect 296646 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 362285 219454
rect 362521 219218 364882 219454
rect 365118 219218 367479 219454
rect 367715 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 434285 219454
rect 434521 219218 436882 219454
rect 437118 219218 439479 219454
rect 439715 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 506285 219454
rect 506521 219218 508882 219454
rect 509118 219218 511479 219454
rect 511715 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 204250 219134
rect 204486 218898 234970 219134
rect 235206 218898 265690 219134
rect 265926 218898 296410 219134
rect 296646 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 362285 219134
rect 362521 218898 364882 219134
rect 365118 218898 367479 219134
rect 367715 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 434285 219134
rect 434521 218898 436882 219134
rect 437118 218898 439479 219134
rect 439715 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 506285 219134
rect 506521 218898 508882 219134
rect 509118 218898 511479 219134
rect 511715 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 219610 201454
rect 219846 201218 250330 201454
rect 250566 201218 281050 201454
rect 281286 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 363583 201454
rect 363819 201218 366180 201454
rect 366416 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 435583 201454
rect 435819 201218 438180 201454
rect 438416 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 507583 201454
rect 507819 201218 510180 201454
rect 510416 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 219610 201134
rect 219846 200898 250330 201134
rect 250566 200898 281050 201134
rect 281286 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 363583 201134
rect 363819 200898 366180 201134
rect 366416 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 435583 201134
rect 435819 200898 438180 201134
rect 438416 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 507583 201134
rect 507819 200898 510180 201134
rect 510416 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 162285 183454
rect 162521 183218 164882 183454
rect 165118 183218 167479 183454
rect 167715 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 204250 183454
rect 204486 183218 234970 183454
rect 235206 183218 265690 183454
rect 265926 183218 296410 183454
rect 296646 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 162285 183134
rect 162521 182898 164882 183134
rect 165118 182898 167479 183134
rect 167715 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 204250 183134
rect 204486 182898 234970 183134
rect 235206 182898 265690 183134
rect 265926 182898 296410 183134
rect 296646 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163583 165454
rect 163819 165218 166180 165454
rect 166416 165218 219610 165454
rect 219846 165218 250330 165454
rect 250566 165218 281050 165454
rect 281286 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163583 165134
rect 163819 164898 166180 165134
rect 166416 164898 219610 165134
rect 219846 164898 250330 165134
rect 250566 164898 281050 165134
rect 281286 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 162285 147454
rect 162521 147218 164882 147454
rect 165118 147218 167479 147454
rect 167715 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 204250 147454
rect 204486 147218 234970 147454
rect 235206 147218 265690 147454
rect 265926 147218 296410 147454
rect 296646 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 362285 147454
rect 362521 147218 364882 147454
rect 365118 147218 367479 147454
rect 367715 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 434285 147454
rect 434521 147218 436882 147454
rect 437118 147218 439479 147454
rect 439715 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 506285 147454
rect 506521 147218 508882 147454
rect 509118 147218 511479 147454
rect 511715 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 162285 147134
rect 162521 146898 164882 147134
rect 165118 146898 167479 147134
rect 167715 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 204250 147134
rect 204486 146898 234970 147134
rect 235206 146898 265690 147134
rect 265926 146898 296410 147134
rect 296646 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 362285 147134
rect 362521 146898 364882 147134
rect 365118 146898 367479 147134
rect 367715 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 434285 147134
rect 434521 146898 436882 147134
rect 437118 146898 439479 147134
rect 439715 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 506285 147134
rect 506521 146898 508882 147134
rect 509118 146898 511479 147134
rect 511715 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163583 129454
rect 163819 129218 166180 129454
rect 166416 129218 219610 129454
rect 219846 129218 250330 129454
rect 250566 129218 281050 129454
rect 281286 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 363583 129454
rect 363819 129218 366180 129454
rect 366416 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 435583 129454
rect 435819 129218 438180 129454
rect 438416 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 507583 129454
rect 507819 129218 510180 129454
rect 510416 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163583 129134
rect 163819 128898 166180 129134
rect 166416 128898 219610 129134
rect 219846 128898 250330 129134
rect 250566 128898 281050 129134
rect 281286 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 363583 129134
rect 363819 128898 366180 129134
rect 366416 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 435583 129134
rect 435819 128898 438180 129134
rect 438416 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 507583 129134
rect 507819 128898 510180 129134
rect 510416 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 204250 111454
rect 204486 111218 234970 111454
rect 235206 111218 265690 111454
rect 265926 111218 296410 111454
rect 296646 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 204250 111134
rect 204486 110898 234970 111134
rect 235206 110898 265690 111134
rect 265926 110898 296410 111134
rect 296646 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use digitalcore_macro  digitalcore
timestamp 1641099986
transform 1 0 200000 0 1 100000
box 0 0 100000 200000
use collapsering_macro  ring0
timestamp 1641099986
transform 1 0 160000 0 1 124000
box 934 0 10000 29776
use ringosc_macro  ring1
timestamp 1641099986
transform 1 0 160000 0 1 160000
box 934 0 10000 29504
use collapsering_macro  ring2
timestamp 1641099986
transform 1 0 360000 0 1 124000
box 934 0 10000 29776
use ringosc_macro  ring3
timestamp 1641099986
transform 1 0 360000 0 1 196000
box 934 0 10000 29504
use collapsering_macro  ring4
timestamp 1641099986
transform 1 0 360000 0 1 268000
box 934 0 10000 29776
use collapsering_macro  ring10
timestamp 1641099986
transform 1 0 432000 0 1 196000
box 934 0 10000 29776
use ringosc_macro  ring11
timestamp 1641099986
transform 1 0 432000 0 1 268000
box 934 0 10000 29504
use ringosc_macro  ring9
timestamp 1641099986
transform 1 0 432000 0 1 124000
box 934 0 10000 29504
use collapsering_macro  ring16
timestamp 1641099986
transform 1 0 504000 0 1 124000
box 934 0 10000 29776
use ringosc_macro  ring17
timestamp 1641099986
transform 1 0 504000 0 1 196000
box 934 0 10000 29504
use collapsering_macro  ring18
timestamp 1641099986
transform 1 0 504000 0 1 268000
box 934 0 10000 29776
use ringosc_macro  ring5
timestamp 1641099986
transform 1 0 360000 0 1 340000
box 934 0 10000 29504
use collapsering_macro  ring6
timestamp 1641099986
transform 1 0 360000 0 1 412000
box 934 0 10000 29776
use ringosc_macro  ring7
timestamp 1641099986
transform 1 0 360000 0 1 484000
box 934 0 10000 29504
use collapsering_macro  ring12
timestamp 1641099986
transform 1 0 432000 0 1 340000
box 934 0 10000 29776
use ringosc_macro  ring13
timestamp 1641099986
transform 1 0 432000 0 1 412000
box 934 0 10000 29504
use collapsering_macro  ring14
timestamp 1641099986
transform 1 0 432000 0 1 484000
box 934 0 10000 29776
use ringosc_macro  ring19
timestamp 1641099986
transform 1 0 504000 0 1 340000
box 934 0 10000 29504
use collapsering_macro  ring20
timestamp 1641099986
transform 1 0 504000 0 1 412000
box 934 0 10000 29776
use ringosc_macro  ring21
timestamp 1641099986
transform 1 0 504000 0 1 484000
box 934 0 10000 29504
use collapsering_macro  ring8
timestamp 1641099986
transform 1 0 360000 0 1 556000
box 934 0 10000 29776
use ringosc_macro  ring15
timestamp 1641099986
transform 1 0 432000 0 1 556000
box 934 0 10000 29504
use collapsering_macro  ring22
timestamp 1641099986
transform 1 0 504000 0 1 556000
box 934 0 10000 29776
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 122000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 156000 362414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 156000 434414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 156000 506414 194000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 228000 362414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 228000 434414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 228000 506414 266000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 300000 362414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 300000 434414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 300000 506414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 372000 362414 410000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 372000 434414 410000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 372000 506414 410000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 444000 362414 482000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 444000 434414 482000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 444000 506414 482000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 516000 362414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 516000 434414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 516000 506414 554000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 302000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 302000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 302000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 588000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 588000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 588000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 122000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 156000 366134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 156000 438134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 156000 510134 194000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 228000 366134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 228000 438134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 228000 510134 266000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 300000 366134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 300000 438134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 300000 510134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 372000 366134 410000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 372000 438134 410000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 372000 510134 410000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 444000 366134 482000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 444000 438134 482000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 444000 510134 482000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 516000 366134 554000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 516000 438134 554000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 516000 510134 554000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 302000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 302000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 302000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 588000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 588000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 588000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 122000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 156000 369854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 156000 441854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 156000 513854 194000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 228000 369854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 228000 441854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 228000 513854 266000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 300000 369854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 300000 441854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 300000 513854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 372000 369854 410000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 372000 441854 410000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 372000 513854 410000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 444000 369854 482000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 444000 441854 482000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 444000 513854 482000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 516000 369854 554000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 516000 441854 554000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 516000 513854 554000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 302000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 302000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 302000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 588000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 588000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 588000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 302000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 302000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 302000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 122000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 156000 171854 158000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 192000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 302000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 302000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 302000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 302000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 302000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 302000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 122000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 156000 164414 158000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 192000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 302000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 302000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 302000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 122000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 156000 168134 158000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 192000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 302000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 302000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 302000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
