magic
tech sky130A
magscale 1 2
timestamp 1641099439
<< obsli1 >>
rect 1104 2159 99147 197489
<< obsm1 >>
rect 106 1300 99898 197520
<< metal2 >>
rect 386 199200 442 200000
rect 1214 199200 1270 200000
rect 2042 199200 2098 200000
rect 2870 199200 2926 200000
rect 3698 199200 3754 200000
rect 4618 199200 4674 200000
rect 5446 199200 5502 200000
rect 6274 199200 6330 200000
rect 7102 199200 7158 200000
rect 7930 199200 7986 200000
rect 8850 199200 8906 200000
rect 9678 199200 9734 200000
rect 10506 199200 10562 200000
rect 11334 199200 11390 200000
rect 12162 199200 12218 200000
rect 13082 199200 13138 200000
rect 13910 199200 13966 200000
rect 14738 199200 14794 200000
rect 15566 199200 15622 200000
rect 16486 199200 16542 200000
rect 17314 199200 17370 200000
rect 18142 199200 18198 200000
rect 18970 199200 19026 200000
rect 19798 199200 19854 200000
rect 20718 199200 20774 200000
rect 21546 199200 21602 200000
rect 22374 199200 22430 200000
rect 23202 199200 23258 200000
rect 24030 199200 24086 200000
rect 24950 199200 25006 200000
rect 25778 199200 25834 200000
rect 26606 199200 26662 200000
rect 27434 199200 27490 200000
rect 28262 199200 28318 200000
rect 29182 199200 29238 200000
rect 30010 199200 30066 200000
rect 30838 199200 30894 200000
rect 31666 199200 31722 200000
rect 32586 199200 32642 200000
rect 33414 199200 33470 200000
rect 34242 199200 34298 200000
rect 35070 199200 35126 200000
rect 35898 199200 35954 200000
rect 36818 199200 36874 200000
rect 37646 199200 37702 200000
rect 38474 199200 38530 200000
rect 39302 199200 39358 200000
rect 40130 199200 40186 200000
rect 41050 199200 41106 200000
rect 41878 199200 41934 200000
rect 42706 199200 42762 200000
rect 43534 199200 43590 200000
rect 44454 199200 44510 200000
rect 45282 199200 45338 200000
rect 46110 199200 46166 200000
rect 46938 199200 46994 200000
rect 47766 199200 47822 200000
rect 48686 199200 48742 200000
rect 49514 199200 49570 200000
rect 50342 199200 50398 200000
rect 51170 199200 51226 200000
rect 51998 199200 52054 200000
rect 52918 199200 52974 200000
rect 53746 199200 53802 200000
rect 54574 199200 54630 200000
rect 55402 199200 55458 200000
rect 56230 199200 56286 200000
rect 57150 199200 57206 200000
rect 57978 199200 58034 200000
rect 58806 199200 58862 200000
rect 59634 199200 59690 200000
rect 60554 199200 60610 200000
rect 61382 199200 61438 200000
rect 62210 199200 62266 200000
rect 63038 199200 63094 200000
rect 63866 199200 63922 200000
rect 64786 199200 64842 200000
rect 65614 199200 65670 200000
rect 66442 199200 66498 200000
rect 67270 199200 67326 200000
rect 68098 199200 68154 200000
rect 69018 199200 69074 200000
rect 69846 199200 69902 200000
rect 70674 199200 70730 200000
rect 71502 199200 71558 200000
rect 72422 199200 72478 200000
rect 73250 199200 73306 200000
rect 74078 199200 74134 200000
rect 74906 199200 74962 200000
rect 75734 199200 75790 200000
rect 76654 199200 76710 200000
rect 77482 199200 77538 200000
rect 78310 199200 78366 200000
rect 79138 199200 79194 200000
rect 79966 199200 80022 200000
rect 80886 199200 80942 200000
rect 81714 199200 81770 200000
rect 82542 199200 82598 200000
rect 83370 199200 83426 200000
rect 84198 199200 84254 200000
rect 85118 199200 85174 200000
rect 85946 199200 86002 200000
rect 86774 199200 86830 200000
rect 87602 199200 87658 200000
rect 88522 199200 88578 200000
rect 89350 199200 89406 200000
rect 90178 199200 90234 200000
rect 91006 199200 91062 200000
rect 91834 199200 91890 200000
rect 92754 199200 92810 200000
rect 93582 199200 93638 200000
rect 94410 199200 94466 200000
rect 95238 199200 95294 200000
rect 96066 199200 96122 200000
rect 96986 199200 97042 200000
rect 97814 199200 97870 200000
rect 98642 199200 98698 200000
rect 99470 199200 99526 200000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7654 0 7710 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18602 0 18658 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64234 0 64290 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81346 0 81402 800
rect 81530 0 81586 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 83922 0 83978 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91466 0 91522 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93490 0 93546 800
rect 93674 0 93730 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95514 0 95570 800
rect 95698 0 95754 800
rect 95882 0 95938 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97906 0 97962 800
rect 98090 0 98146 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 199144 330 199200
rect 498 199144 1158 199200
rect 1326 199144 1986 199200
rect 2154 199144 2814 199200
rect 2982 199144 3642 199200
rect 3810 199144 4562 199200
rect 4730 199144 5390 199200
rect 5558 199144 6218 199200
rect 6386 199144 7046 199200
rect 7214 199144 7874 199200
rect 8042 199144 8794 199200
rect 8962 199144 9622 199200
rect 9790 199144 10450 199200
rect 10618 199144 11278 199200
rect 11446 199144 12106 199200
rect 12274 199144 13026 199200
rect 13194 199144 13854 199200
rect 14022 199144 14682 199200
rect 14850 199144 15510 199200
rect 15678 199144 16430 199200
rect 16598 199144 17258 199200
rect 17426 199144 18086 199200
rect 18254 199144 18914 199200
rect 19082 199144 19742 199200
rect 19910 199144 20662 199200
rect 20830 199144 21490 199200
rect 21658 199144 22318 199200
rect 22486 199144 23146 199200
rect 23314 199144 23974 199200
rect 24142 199144 24894 199200
rect 25062 199144 25722 199200
rect 25890 199144 26550 199200
rect 26718 199144 27378 199200
rect 27546 199144 28206 199200
rect 28374 199144 29126 199200
rect 29294 199144 29954 199200
rect 30122 199144 30782 199200
rect 30950 199144 31610 199200
rect 31778 199144 32530 199200
rect 32698 199144 33358 199200
rect 33526 199144 34186 199200
rect 34354 199144 35014 199200
rect 35182 199144 35842 199200
rect 36010 199144 36762 199200
rect 36930 199144 37590 199200
rect 37758 199144 38418 199200
rect 38586 199144 39246 199200
rect 39414 199144 40074 199200
rect 40242 199144 40994 199200
rect 41162 199144 41822 199200
rect 41990 199144 42650 199200
rect 42818 199144 43478 199200
rect 43646 199144 44398 199200
rect 44566 199144 45226 199200
rect 45394 199144 46054 199200
rect 46222 199144 46882 199200
rect 47050 199144 47710 199200
rect 47878 199144 48630 199200
rect 48798 199144 49458 199200
rect 49626 199144 50286 199200
rect 50454 199144 51114 199200
rect 51282 199144 51942 199200
rect 52110 199144 52862 199200
rect 53030 199144 53690 199200
rect 53858 199144 54518 199200
rect 54686 199144 55346 199200
rect 55514 199144 56174 199200
rect 56342 199144 57094 199200
rect 57262 199144 57922 199200
rect 58090 199144 58750 199200
rect 58918 199144 59578 199200
rect 59746 199144 60498 199200
rect 60666 199144 61326 199200
rect 61494 199144 62154 199200
rect 62322 199144 62982 199200
rect 63150 199144 63810 199200
rect 63978 199144 64730 199200
rect 64898 199144 65558 199200
rect 65726 199144 66386 199200
rect 66554 199144 67214 199200
rect 67382 199144 68042 199200
rect 68210 199144 68962 199200
rect 69130 199144 69790 199200
rect 69958 199144 70618 199200
rect 70786 199144 71446 199200
rect 71614 199144 72366 199200
rect 72534 199144 73194 199200
rect 73362 199144 74022 199200
rect 74190 199144 74850 199200
rect 75018 199144 75678 199200
rect 75846 199144 76598 199200
rect 76766 199144 77426 199200
rect 77594 199144 78254 199200
rect 78422 199144 79082 199200
rect 79250 199144 79910 199200
rect 80078 199144 80830 199200
rect 80998 199144 81658 199200
rect 81826 199144 82486 199200
rect 82654 199144 83314 199200
rect 83482 199144 84142 199200
rect 84310 199144 85062 199200
rect 85230 199144 85890 199200
rect 86058 199144 86718 199200
rect 86886 199144 87546 199200
rect 87714 199144 88466 199200
rect 88634 199144 89294 199200
rect 89462 199144 90122 199200
rect 90290 199144 90950 199200
rect 91118 199144 91778 199200
rect 91946 199144 92698 199200
rect 92866 199144 93526 199200
rect 93694 199144 94354 199200
rect 94522 199144 95182 199200
rect 95350 199144 96010 199200
rect 96178 199144 96930 199200
rect 97098 199144 97758 199200
rect 97926 199144 98586 199200
rect 98754 199144 99414 199200
rect 99582 199144 99892 199200
rect 112 856 99892 199144
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 974 856
rect 1142 800 1158 856
rect 1326 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 1986 856
rect 2154 800 2170 856
rect 2338 800 2354 856
rect 2522 800 2630 856
rect 2798 800 2814 856
rect 2982 800 2998 856
rect 3166 800 3182 856
rect 3350 800 3366 856
rect 3534 800 3550 856
rect 3718 800 3826 856
rect 3994 800 4010 856
rect 4178 800 4194 856
rect 4362 800 4378 856
rect 4546 800 4562 856
rect 4730 800 4746 856
rect 4914 800 5022 856
rect 5190 800 5206 856
rect 5374 800 5390 856
rect 5558 800 5574 856
rect 5742 800 5758 856
rect 5926 800 5942 856
rect 6110 800 6218 856
rect 6386 800 6402 856
rect 6570 800 6586 856
rect 6754 800 6770 856
rect 6938 800 6954 856
rect 7122 800 7138 856
rect 7306 800 7414 856
rect 7582 800 7598 856
rect 7766 800 7782 856
rect 7950 800 7966 856
rect 8134 800 8150 856
rect 8318 800 8334 856
rect 8502 800 8610 856
rect 8778 800 8794 856
rect 8962 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9530 856
rect 9698 800 9806 856
rect 9974 800 9990 856
rect 10158 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10726 856
rect 10894 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11554 856
rect 11722 800 11738 856
rect 11906 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12566 856
rect 12734 800 12750 856
rect 12918 800 12934 856
rect 13102 800 13118 856
rect 13286 800 13394 856
rect 13562 800 13578 856
rect 13746 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14130 856
rect 14298 800 14314 856
rect 14482 800 14590 856
rect 14758 800 14774 856
rect 14942 800 14958 856
rect 15126 800 15142 856
rect 15310 800 15326 856
rect 15494 800 15510 856
rect 15678 800 15786 856
rect 15954 800 15970 856
rect 16138 800 16154 856
rect 16322 800 16338 856
rect 16506 800 16522 856
rect 16690 800 16706 856
rect 16874 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17350 856
rect 17518 800 17534 856
rect 17702 800 17718 856
rect 17886 800 17902 856
rect 18070 800 18178 856
rect 18346 800 18362 856
rect 18530 800 18546 856
rect 18714 800 18730 856
rect 18898 800 18914 856
rect 19082 800 19098 856
rect 19266 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20110 856
rect 20278 800 20294 856
rect 20462 800 20570 856
rect 20738 800 20754 856
rect 20922 800 20938 856
rect 21106 800 21122 856
rect 21290 800 21306 856
rect 21474 800 21490 856
rect 21658 800 21766 856
rect 21934 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22318 856
rect 22486 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22962 856
rect 23130 800 23146 856
rect 23314 800 23330 856
rect 23498 800 23514 856
rect 23682 800 23698 856
rect 23866 800 23882 856
rect 24050 800 24158 856
rect 24326 800 24342 856
rect 24510 800 24526 856
rect 24694 800 24710 856
rect 24878 800 24894 856
rect 25062 800 25078 856
rect 25246 800 25262 856
rect 25430 800 25538 856
rect 25706 800 25722 856
rect 25890 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26274 856
rect 26442 800 26458 856
rect 26626 800 26734 856
rect 26902 800 26918 856
rect 27086 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28666 856
rect 28834 800 28850 856
rect 29018 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29494 856
rect 29662 800 29678 856
rect 29846 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30322 856
rect 30490 800 30506 856
rect 30674 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31058 856
rect 31226 800 31242 856
rect 31410 800 31518 856
rect 31686 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32070 856
rect 32238 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32714 856
rect 32882 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33266 856
rect 33434 800 33450 856
rect 33618 800 33634 856
rect 33802 800 33910 856
rect 34078 800 34094 856
rect 34262 800 34278 856
rect 34446 800 34462 856
rect 34630 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35106 856
rect 35274 800 35290 856
rect 35458 800 35474 856
rect 35642 800 35658 856
rect 35826 800 35842 856
rect 36010 800 36026 856
rect 36194 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36854 856
rect 37022 800 37038 856
rect 37206 800 37222 856
rect 37390 800 37498 856
rect 37666 800 37682 856
rect 37850 800 37866 856
rect 38034 800 38050 856
rect 38218 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39062 856
rect 39230 800 39246 856
rect 39414 800 39430 856
rect 39598 800 39614 856
rect 39782 800 39890 856
rect 40058 800 40074 856
rect 40242 800 40258 856
rect 40426 800 40442 856
rect 40610 800 40626 856
rect 40794 800 40810 856
rect 40978 800 41086 856
rect 41254 800 41270 856
rect 41438 800 41454 856
rect 41622 800 41638 856
rect 41806 800 41822 856
rect 41990 800 42006 856
rect 42174 800 42282 856
rect 42450 800 42466 856
rect 42634 800 42650 856
rect 42818 800 42834 856
rect 43002 800 43018 856
rect 43186 800 43202 856
rect 43370 800 43478 856
rect 43646 800 43662 856
rect 43830 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44398 856
rect 44566 800 44674 856
rect 44842 800 44858 856
rect 45026 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45410 856
rect 45578 800 45594 856
rect 45762 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46238 856
rect 46406 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46790 856
rect 46958 800 47066 856
rect 47234 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47618 856
rect 47786 800 47802 856
rect 47970 800 47986 856
rect 48154 800 48262 856
rect 48430 800 48446 856
rect 48614 800 48630 856
rect 48798 800 48814 856
rect 48982 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49458 856
rect 49626 800 49642 856
rect 49810 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50194 856
rect 50362 800 50378 856
rect 50546 800 50562 856
rect 50730 800 50838 856
rect 51006 800 51022 856
rect 51190 800 51206 856
rect 51374 800 51390 856
rect 51558 800 51574 856
rect 51742 800 51758 856
rect 51926 800 52034 856
rect 52202 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52586 856
rect 52754 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53230 856
rect 53398 800 53414 856
rect 53582 800 53598 856
rect 53766 800 53782 856
rect 53950 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54426 856
rect 54594 800 54610 856
rect 54778 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55162 856
rect 55330 800 55346 856
rect 55514 800 55622 856
rect 55790 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56174 856
rect 56342 800 56358 856
rect 56526 800 56542 856
rect 56710 800 56818 856
rect 56986 800 57002 856
rect 57170 800 57186 856
rect 57354 800 57370 856
rect 57538 800 57554 856
rect 57722 800 57738 856
rect 57906 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58382 856
rect 58550 800 58566 856
rect 58734 800 58750 856
rect 58918 800 58934 856
rect 59102 800 59210 856
rect 59378 800 59394 856
rect 59562 800 59578 856
rect 59746 800 59762 856
rect 59930 800 59946 856
rect 60114 800 60130 856
rect 60298 800 60406 856
rect 60574 800 60590 856
rect 60758 800 60774 856
rect 60942 800 60958 856
rect 61126 800 61142 856
rect 61310 800 61326 856
rect 61494 800 61602 856
rect 61770 800 61786 856
rect 61954 800 61970 856
rect 62138 800 62154 856
rect 62322 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62798 856
rect 62966 800 62982 856
rect 63150 800 63166 856
rect 63334 800 63350 856
rect 63518 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63994 856
rect 64162 800 64178 856
rect 64346 800 64362 856
rect 64530 800 64546 856
rect 64714 800 64730 856
rect 64898 800 64914 856
rect 65082 800 65190 856
rect 65358 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66110 856
rect 66278 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66754 856
rect 66922 800 66938 856
rect 67106 800 67122 856
rect 67290 800 67306 856
rect 67474 800 67582 856
rect 67750 800 67766 856
rect 67934 800 67950 856
rect 68118 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68778 856
rect 68946 800 68962 856
rect 69130 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69514 856
rect 69682 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70342 856
rect 70510 800 70526 856
rect 70694 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71170 856
rect 71338 800 71354 856
rect 71522 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71906 856
rect 72074 800 72090 856
rect 72258 800 72366 856
rect 72534 800 72550 856
rect 72718 800 72734 856
rect 72902 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73286 856
rect 73454 800 73562 856
rect 73730 800 73746 856
rect 73914 800 73930 856
rect 74098 800 74114 856
rect 74282 800 74298 856
rect 74466 800 74482 856
rect 74650 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75310 856
rect 75478 800 75494 856
rect 75662 800 75678 856
rect 75846 800 75862 856
rect 76030 800 76138 856
rect 76306 800 76322 856
rect 76490 800 76506 856
rect 76674 800 76690 856
rect 76858 800 76874 856
rect 77042 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77518 856
rect 77686 800 77702 856
rect 77870 800 77886 856
rect 78054 800 78070 856
rect 78238 800 78254 856
rect 78422 800 78530 856
rect 78698 800 78714 856
rect 78882 800 78898 856
rect 79066 800 79082 856
rect 79250 800 79266 856
rect 79434 800 79450 856
rect 79618 800 79726 856
rect 79894 800 79910 856
rect 80078 800 80094 856
rect 80262 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80646 856
rect 80814 800 80922 856
rect 81090 800 81106 856
rect 81274 800 81290 856
rect 81458 800 81474 856
rect 81642 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82118 856
rect 82286 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82854 856
rect 83022 800 83038 856
rect 83206 800 83314 856
rect 83482 800 83498 856
rect 83666 800 83682 856
rect 83850 800 83866 856
rect 84034 800 84050 856
rect 84218 800 84234 856
rect 84402 800 84510 856
rect 84678 800 84694 856
rect 84862 800 84878 856
rect 85046 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85430 856
rect 85598 800 85706 856
rect 85874 800 85890 856
rect 86058 800 86074 856
rect 86242 800 86258 856
rect 86426 800 86442 856
rect 86610 800 86626 856
rect 86794 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88098 856
rect 88266 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88650 856
rect 88818 800 88834 856
rect 89002 800 89018 856
rect 89186 800 89294 856
rect 89462 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90214 856
rect 90382 800 90490 856
rect 90658 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91042 856
rect 91210 800 91226 856
rect 91394 800 91410 856
rect 91578 800 91686 856
rect 91854 800 91870 856
rect 92038 800 92054 856
rect 92222 800 92238 856
rect 92406 800 92422 856
rect 92590 800 92606 856
rect 92774 800 92882 856
rect 93050 800 93066 856
rect 93234 800 93250 856
rect 93418 800 93434 856
rect 93602 800 93618 856
rect 93786 800 93802 856
rect 93970 800 94078 856
rect 94246 800 94262 856
rect 94430 800 94446 856
rect 94614 800 94630 856
rect 94798 800 94814 856
rect 94982 800 94998 856
rect 95166 800 95274 856
rect 95442 800 95458 856
rect 95626 800 95642 856
rect 95810 800 95826 856
rect 95994 800 96010 856
rect 96178 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96654 856
rect 96822 800 96838 856
rect 97006 800 97022 856
rect 97190 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97666 856
rect 97834 800 97850 856
rect 98018 800 98034 856
rect 98202 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98862 856
rect 99030 800 99046 856
rect 99214 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 198840 800 198960
rect 99200 198432 100000 198552
rect 0 196800 800 196920
rect 99200 195304 100000 195424
rect 0 194624 800 194744
rect 0 192584 800 192704
rect 99200 192312 100000 192432
rect 0 190408 800 190528
rect 99200 189184 100000 189304
rect 0 188368 800 188488
rect 0 186192 800 186312
rect 99200 186056 100000 186176
rect 0 184152 800 184272
rect 99200 183064 100000 183184
rect 0 181976 800 182096
rect 0 179936 800 180056
rect 99200 179936 100000 180056
rect 0 177760 800 177880
rect 99200 176808 100000 176928
rect 0 175720 800 175840
rect 99200 173816 100000 173936
rect 0 173544 800 173664
rect 0 171504 800 171624
rect 99200 170688 100000 170808
rect 0 169328 800 169448
rect 99200 167696 100000 167816
rect 0 167288 800 167408
rect 0 165112 800 165232
rect 99200 164568 100000 164688
rect 0 163072 800 163192
rect 99200 161440 100000 161560
rect 0 160896 800 161016
rect 0 158856 800 158976
rect 99200 158448 100000 158568
rect 0 156680 800 156800
rect 99200 155320 100000 155440
rect 0 154640 800 154760
rect 0 152464 800 152584
rect 99200 152192 100000 152312
rect 0 150424 800 150544
rect 99200 149200 100000 149320
rect 0 148248 800 148368
rect 0 146208 800 146328
rect 99200 146072 100000 146192
rect 0 144032 800 144152
rect 99200 143080 100000 143200
rect 0 141992 800 142112
rect 0 139816 800 139936
rect 99200 139952 100000 140072
rect 0 137776 800 137896
rect 99200 136824 100000 136944
rect 0 135600 800 135720
rect 99200 133832 100000 133952
rect 0 133560 800 133680
rect 0 131520 800 131640
rect 99200 130704 100000 130824
rect 0 129344 800 129464
rect 99200 127576 100000 127696
rect 0 127304 800 127424
rect 0 125128 800 125248
rect 99200 124584 100000 124704
rect 0 123088 800 123208
rect 99200 121456 100000 121576
rect 0 120912 800 121032
rect 0 118872 800 118992
rect 99200 118328 100000 118448
rect 0 116696 800 116816
rect 99200 115336 100000 115456
rect 0 114656 800 114776
rect 0 112480 800 112600
rect 99200 112208 100000 112328
rect 0 110440 800 110560
rect 99200 109216 100000 109336
rect 0 108264 800 108384
rect 0 106224 800 106344
rect 99200 106088 100000 106208
rect 0 104048 800 104168
rect 99200 102960 100000 103080
rect 0 102008 800 102128
rect 0 99832 800 99952
rect 99200 99968 100000 100088
rect 0 97792 800 97912
rect 99200 96840 100000 96960
rect 0 95616 800 95736
rect 0 93576 800 93696
rect 99200 93712 100000 93832
rect 0 91400 800 91520
rect 99200 90720 100000 90840
rect 0 89360 800 89480
rect 99200 87592 100000 87712
rect 0 87184 800 87304
rect 0 85144 800 85264
rect 99200 84600 100000 84720
rect 0 82968 800 83088
rect 99200 81472 100000 81592
rect 0 80928 800 81048
rect 0 78752 800 78872
rect 99200 78344 100000 78464
rect 0 76712 800 76832
rect 99200 75352 100000 75472
rect 0 74536 800 74656
rect 0 72496 800 72616
rect 99200 72224 100000 72344
rect 0 70320 800 70440
rect 99200 69096 100000 69216
rect 0 68280 800 68400
rect 0 66240 800 66360
rect 99200 66104 100000 66224
rect 0 64064 800 64184
rect 99200 62976 100000 63096
rect 0 62024 800 62144
rect 0 59848 800 59968
rect 99200 59848 100000 59968
rect 0 57808 800 57928
rect 99200 56856 100000 56976
rect 0 55632 800 55752
rect 0 53592 800 53712
rect 99200 53728 100000 53848
rect 0 51416 800 51536
rect 99200 50736 100000 50856
rect 0 49376 800 49496
rect 99200 47608 100000 47728
rect 0 47200 800 47320
rect 0 45160 800 45280
rect 99200 44480 100000 44600
rect 0 42984 800 43104
rect 99200 41488 100000 41608
rect 0 40944 800 41064
rect 0 38768 800 38888
rect 99200 38360 100000 38480
rect 0 36728 800 36848
rect 99200 35232 100000 35352
rect 0 34552 800 34672
rect 0 32512 800 32632
rect 99200 32240 100000 32360
rect 0 30336 800 30456
rect 99200 29112 100000 29232
rect 0 28296 800 28416
rect 0 26120 800 26240
rect 99200 26120 100000 26240
rect 0 24080 800 24200
rect 99200 22992 100000 23112
rect 0 21904 800 22024
rect 0 19864 800 19984
rect 99200 19864 100000 19984
rect 0 17688 800 17808
rect 99200 16872 100000 16992
rect 0 15648 800 15768
rect 99200 13744 100000 13864
rect 0 13472 800 13592
rect 0 11432 800 11552
rect 99200 10616 100000 10736
rect 0 9256 800 9376
rect 99200 7624 100000 7744
rect 0 7216 800 7336
rect 0 5040 800 5160
rect 99200 4496 100000 4616
rect 0 3000 800 3120
rect 99200 1504 100000 1624
rect 0 960 800 1080
<< obsm3 >>
rect 880 198760 99200 198933
rect 798 198632 99200 198760
rect 798 198352 99120 198632
rect 798 197000 99200 198352
rect 880 196720 99200 197000
rect 798 195504 99200 196720
rect 798 195224 99120 195504
rect 798 194824 99200 195224
rect 880 194544 99200 194824
rect 798 192784 99200 194544
rect 880 192512 99200 192784
rect 880 192504 99120 192512
rect 798 192232 99120 192504
rect 798 190608 99200 192232
rect 880 190328 99200 190608
rect 798 189384 99200 190328
rect 798 189104 99120 189384
rect 798 188568 99200 189104
rect 880 188288 99200 188568
rect 798 186392 99200 188288
rect 880 186256 99200 186392
rect 880 186112 99120 186256
rect 798 185976 99120 186112
rect 798 184352 99200 185976
rect 880 184072 99200 184352
rect 798 183264 99200 184072
rect 798 182984 99120 183264
rect 798 182176 99200 182984
rect 880 181896 99200 182176
rect 798 180136 99200 181896
rect 880 179856 99120 180136
rect 798 177960 99200 179856
rect 880 177680 99200 177960
rect 798 177008 99200 177680
rect 798 176728 99120 177008
rect 798 175920 99200 176728
rect 880 175640 99200 175920
rect 798 174016 99200 175640
rect 798 173744 99120 174016
rect 880 173736 99120 173744
rect 880 173464 99200 173736
rect 798 171704 99200 173464
rect 880 171424 99200 171704
rect 798 170888 99200 171424
rect 798 170608 99120 170888
rect 798 169528 99200 170608
rect 880 169248 99200 169528
rect 798 167896 99200 169248
rect 798 167616 99120 167896
rect 798 167488 99200 167616
rect 880 167208 99200 167488
rect 798 165312 99200 167208
rect 880 165032 99200 165312
rect 798 164768 99200 165032
rect 798 164488 99120 164768
rect 798 163272 99200 164488
rect 880 162992 99200 163272
rect 798 161640 99200 162992
rect 798 161360 99120 161640
rect 798 161096 99200 161360
rect 880 160816 99200 161096
rect 798 159056 99200 160816
rect 880 158776 99200 159056
rect 798 158648 99200 158776
rect 798 158368 99120 158648
rect 798 156880 99200 158368
rect 880 156600 99200 156880
rect 798 155520 99200 156600
rect 798 155240 99120 155520
rect 798 154840 99200 155240
rect 880 154560 99200 154840
rect 798 152664 99200 154560
rect 880 152392 99200 152664
rect 880 152384 99120 152392
rect 798 152112 99120 152384
rect 798 150624 99200 152112
rect 880 150344 99200 150624
rect 798 149400 99200 150344
rect 798 149120 99120 149400
rect 798 148448 99200 149120
rect 880 148168 99200 148448
rect 798 146408 99200 148168
rect 880 146272 99200 146408
rect 880 146128 99120 146272
rect 798 145992 99120 146128
rect 798 144232 99200 145992
rect 880 143952 99200 144232
rect 798 143280 99200 143952
rect 798 143000 99120 143280
rect 798 142192 99200 143000
rect 880 141912 99200 142192
rect 798 140152 99200 141912
rect 798 140016 99120 140152
rect 880 139872 99120 140016
rect 880 139736 99200 139872
rect 798 137976 99200 139736
rect 880 137696 99200 137976
rect 798 137024 99200 137696
rect 798 136744 99120 137024
rect 798 135800 99200 136744
rect 880 135520 99200 135800
rect 798 134032 99200 135520
rect 798 133760 99120 134032
rect 880 133752 99120 133760
rect 880 133480 99200 133752
rect 798 131720 99200 133480
rect 880 131440 99200 131720
rect 798 130904 99200 131440
rect 798 130624 99120 130904
rect 798 129544 99200 130624
rect 880 129264 99200 129544
rect 798 127776 99200 129264
rect 798 127504 99120 127776
rect 880 127496 99120 127504
rect 880 127224 99200 127496
rect 798 125328 99200 127224
rect 880 125048 99200 125328
rect 798 124784 99200 125048
rect 798 124504 99120 124784
rect 798 123288 99200 124504
rect 880 123008 99200 123288
rect 798 121656 99200 123008
rect 798 121376 99120 121656
rect 798 121112 99200 121376
rect 880 120832 99200 121112
rect 798 119072 99200 120832
rect 880 118792 99200 119072
rect 798 118528 99200 118792
rect 798 118248 99120 118528
rect 798 116896 99200 118248
rect 880 116616 99200 116896
rect 798 115536 99200 116616
rect 798 115256 99120 115536
rect 798 114856 99200 115256
rect 880 114576 99200 114856
rect 798 112680 99200 114576
rect 880 112408 99200 112680
rect 880 112400 99120 112408
rect 798 112128 99120 112400
rect 798 110640 99200 112128
rect 880 110360 99200 110640
rect 798 109416 99200 110360
rect 798 109136 99120 109416
rect 798 108464 99200 109136
rect 880 108184 99200 108464
rect 798 106424 99200 108184
rect 880 106288 99200 106424
rect 880 106144 99120 106288
rect 798 106008 99120 106144
rect 798 104248 99200 106008
rect 880 103968 99200 104248
rect 798 103160 99200 103968
rect 798 102880 99120 103160
rect 798 102208 99200 102880
rect 880 101928 99200 102208
rect 798 100168 99200 101928
rect 798 100032 99120 100168
rect 880 99888 99120 100032
rect 880 99752 99200 99888
rect 798 97992 99200 99752
rect 880 97712 99200 97992
rect 798 97040 99200 97712
rect 798 96760 99120 97040
rect 798 95816 99200 96760
rect 880 95536 99200 95816
rect 798 93912 99200 95536
rect 798 93776 99120 93912
rect 880 93632 99120 93776
rect 880 93496 99200 93632
rect 798 91600 99200 93496
rect 880 91320 99200 91600
rect 798 90920 99200 91320
rect 798 90640 99120 90920
rect 798 89560 99200 90640
rect 880 89280 99200 89560
rect 798 87792 99200 89280
rect 798 87512 99120 87792
rect 798 87384 99200 87512
rect 880 87104 99200 87384
rect 798 85344 99200 87104
rect 880 85064 99200 85344
rect 798 84800 99200 85064
rect 798 84520 99120 84800
rect 798 83168 99200 84520
rect 880 82888 99200 83168
rect 798 81672 99200 82888
rect 798 81392 99120 81672
rect 798 81128 99200 81392
rect 880 80848 99200 81128
rect 798 78952 99200 80848
rect 880 78672 99200 78952
rect 798 78544 99200 78672
rect 798 78264 99120 78544
rect 798 76912 99200 78264
rect 880 76632 99200 76912
rect 798 75552 99200 76632
rect 798 75272 99120 75552
rect 798 74736 99200 75272
rect 880 74456 99200 74736
rect 798 72696 99200 74456
rect 880 72424 99200 72696
rect 880 72416 99120 72424
rect 798 72144 99120 72416
rect 798 70520 99200 72144
rect 880 70240 99200 70520
rect 798 69296 99200 70240
rect 798 69016 99120 69296
rect 798 68480 99200 69016
rect 880 68200 99200 68480
rect 798 66440 99200 68200
rect 880 66304 99200 66440
rect 880 66160 99120 66304
rect 798 66024 99120 66160
rect 798 64264 99200 66024
rect 880 63984 99200 64264
rect 798 63176 99200 63984
rect 798 62896 99120 63176
rect 798 62224 99200 62896
rect 880 61944 99200 62224
rect 798 60048 99200 61944
rect 880 59768 99120 60048
rect 798 58008 99200 59768
rect 880 57728 99200 58008
rect 798 57056 99200 57728
rect 798 56776 99120 57056
rect 798 55832 99200 56776
rect 880 55552 99200 55832
rect 798 53928 99200 55552
rect 798 53792 99120 53928
rect 880 53648 99120 53792
rect 880 53512 99200 53648
rect 798 51616 99200 53512
rect 880 51336 99200 51616
rect 798 50936 99200 51336
rect 798 50656 99120 50936
rect 798 49576 99200 50656
rect 880 49296 99200 49576
rect 798 47808 99200 49296
rect 798 47528 99120 47808
rect 798 47400 99200 47528
rect 880 47120 99200 47400
rect 798 45360 99200 47120
rect 880 45080 99200 45360
rect 798 44680 99200 45080
rect 798 44400 99120 44680
rect 798 43184 99200 44400
rect 880 42904 99200 43184
rect 798 41688 99200 42904
rect 798 41408 99120 41688
rect 798 41144 99200 41408
rect 880 40864 99200 41144
rect 798 38968 99200 40864
rect 880 38688 99200 38968
rect 798 38560 99200 38688
rect 798 38280 99120 38560
rect 798 36928 99200 38280
rect 880 36648 99200 36928
rect 798 35432 99200 36648
rect 798 35152 99120 35432
rect 798 34752 99200 35152
rect 880 34472 99200 34752
rect 798 32712 99200 34472
rect 880 32440 99200 32712
rect 880 32432 99120 32440
rect 798 32160 99120 32432
rect 798 30536 99200 32160
rect 880 30256 99200 30536
rect 798 29312 99200 30256
rect 798 29032 99120 29312
rect 798 28496 99200 29032
rect 880 28216 99200 28496
rect 798 26320 99200 28216
rect 880 26040 99120 26320
rect 798 24280 99200 26040
rect 880 24000 99200 24280
rect 798 23192 99200 24000
rect 798 22912 99120 23192
rect 798 22104 99200 22912
rect 880 21824 99200 22104
rect 798 20064 99200 21824
rect 880 19784 99120 20064
rect 798 17888 99200 19784
rect 880 17608 99200 17888
rect 798 17072 99200 17608
rect 798 16792 99120 17072
rect 798 15848 99200 16792
rect 880 15568 99200 15848
rect 798 13944 99200 15568
rect 798 13672 99120 13944
rect 880 13664 99120 13672
rect 880 13392 99200 13664
rect 798 11632 99200 13392
rect 880 11352 99200 11632
rect 798 10816 99200 11352
rect 798 10536 99120 10816
rect 798 9456 99200 10536
rect 880 9176 99200 9456
rect 798 7824 99200 9176
rect 798 7544 99120 7824
rect 798 7416 99200 7544
rect 880 7136 99200 7416
rect 798 5240 99200 7136
rect 880 4960 99200 5240
rect 798 4696 99200 4960
rect 798 4416 99120 4696
rect 798 3200 99200 4416
rect 880 2920 99200 3200
rect 798 1704 99200 2920
rect 798 1424 99120 1704
rect 798 1160 99200 1424
rect 880 987 99200 1160
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
<< obsm4 >>
rect 1715 2347 4128 191589
rect 4608 2347 19488 191589
rect 19968 2347 34848 191589
rect 35328 2347 50208 191589
rect 50688 2347 65568 191589
rect 66048 2347 80928 191589
rect 81408 2347 96173 191589
<< labels >>
rlabel metal2 s 386 199200 442 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 25778 199200 25834 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 28262 199200 28318 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 30838 199200 30894 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 33414 199200 33470 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 35898 199200 35954 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 38474 199200 38530 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 41050 199200 41106 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 43534 199200 43590 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 46110 199200 46166 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 48686 199200 48742 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2870 199200 2926 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 51170 199200 51226 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 53746 199200 53802 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 56230 199200 56286 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 58806 199200 58862 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 61382 199200 61438 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 63866 199200 63922 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 66442 199200 66498 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 69018 199200 69074 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 71502 199200 71558 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 74078 199200 74134 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5446 199200 5502 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 76654 199200 76710 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 79138 199200 79194 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 81714 199200 81770 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 84198 199200 84254 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 86774 199200 86830 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 89350 199200 89406 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 91834 199200 91890 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 94410 199200 94466 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7930 199200 7986 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10506 199200 10562 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13082 199200 13138 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 15566 199200 15622 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18142 199200 18198 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 20718 199200 20774 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23202 199200 23258 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 199200 1270 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 26606 199200 26662 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 29182 199200 29238 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 31666 199200 31722 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 34242 199200 34298 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 36818 199200 36874 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 39302 199200 39358 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 41878 199200 41934 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 44454 199200 44510 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 46938 199200 46994 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 49514 199200 49570 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3698 199200 3754 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 51998 199200 52054 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 54574 199200 54630 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 57150 199200 57206 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 59634 199200 59690 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 62210 199200 62266 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 64786 199200 64842 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 67270 199200 67326 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 69846 199200 69902 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 72422 199200 72478 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 74906 199200 74962 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6274 199200 6330 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 77482 199200 77538 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 79966 199200 80022 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 82542 199200 82598 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 85118 199200 85174 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 87602 199200 87658 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 90178 199200 90234 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 92754 199200 92810 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 95238 199200 95294 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8850 199200 8906 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11334 199200 11390 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13910 199200 13966 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 16486 199200 16542 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 18970 199200 19026 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 21546 199200 21602 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24030 199200 24086 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2042 199200 2098 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 27434 199200 27490 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 30010 199200 30066 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 32586 199200 32642 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 35070 199200 35126 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 37646 199200 37702 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 40130 199200 40186 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 42706 199200 42762 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 45282 199200 45338 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 47766 199200 47822 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 50342 199200 50398 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4618 199200 4674 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 52918 199200 52974 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 55402 199200 55458 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 57978 199200 58034 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 60554 199200 60610 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 63038 199200 63094 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 65614 199200 65670 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 68098 199200 68154 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 70674 199200 70730 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 73250 199200 73306 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 75734 199200 75790 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7102 199200 7158 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 78310 199200 78366 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 80886 199200 80942 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 83370 199200 83426 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 85946 199200 86002 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 88522 199200 88578 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 91006 199200 91062 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 93582 199200 93638 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 96066 199200 96122 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9678 199200 9734 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12162 199200 12218 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14738 199200 14794 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17314 199200 17370 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 19798 199200 19854 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22374 199200 22430 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 24950 199200 25006 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 ring0_clk
port 502 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 ring0_clkmux[0]
port 503 nsew signal output
rlabel metal3 s 0 120912 800 121032 6 ring0_clkmux[1]
port 504 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 ring0_clkmux[2]
port 505 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 ring0_start
port 506 nsew signal output
rlabel metal3 s 0 960 800 1080 6 ring0_trim_a[0]
port 507 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 ring0_trim_a[10]
port 508 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 ring0_trim_a[11]
port 509 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 ring0_trim_a[12]
port 510 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 ring0_trim_a[13]
port 511 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 ring0_trim_a[14]
port 512 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 ring0_trim_a[15]
port 513 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 ring0_trim_a[16]
port 514 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 ring0_trim_a[17]
port 515 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 ring0_trim_a[18]
port 516 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 ring0_trim_a[19]
port 517 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 ring0_trim_a[1]
port 518 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 ring0_trim_a[20]
port 519 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 ring0_trim_a[21]
port 520 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 ring0_trim_a[22]
port 521 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 ring0_trim_a[23]
port 522 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 ring0_trim_a[24]
port 523 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 ring0_trim_a[25]
port 524 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 ring0_trim_a[26]
port 525 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 ring0_trim_a[27]
port 526 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 ring0_trim_a[2]
port 527 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 ring0_trim_a[3]
port 528 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 ring0_trim_a[4]
port 529 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 ring0_trim_a[5]
port 530 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 ring0_trim_a[6]
port 531 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 ring0_trim_a[7]
port 532 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 ring0_trim_a[8]
port 533 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 ring0_trim_a[9]
port 534 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 ring0_trim_b[0]
port 535 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 ring0_trim_b[10]
port 536 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 ring0_trim_b[11]
port 537 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 ring0_trim_b[12]
port 538 nsew signal output
rlabel metal3 s 0 87184 800 87304 6 ring0_trim_b[13]
port 539 nsew signal output
rlabel metal3 s 0 89360 800 89480 6 ring0_trim_b[14]
port 540 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 ring0_trim_b[15]
port 541 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 ring0_trim_b[16]
port 542 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 ring0_trim_b[17]
port 543 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 ring0_trim_b[18]
port 544 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 ring0_trim_b[19]
port 545 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 ring0_trim_b[1]
port 546 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 ring0_trim_b[20]
port 547 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 ring0_trim_b[21]
port 548 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 ring0_trim_b[22]
port 549 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 ring0_trim_b[23]
port 550 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 ring0_trim_b[24]
port 551 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 ring0_trim_b[25]
port 552 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 ring0_trim_b[26]
port 553 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 ring0_trim_b[27]
port 554 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 ring0_trim_b[2]
port 555 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 ring0_trim_b[3]
port 556 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 ring0_trim_b[4]
port 557 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 ring0_trim_b[5]
port 558 nsew signal output
rlabel metal3 s 0 72496 800 72616 6 ring0_trim_b[6]
port 559 nsew signal output
rlabel metal3 s 0 74536 800 74656 6 ring0_trim_b[7]
port 560 nsew signal output
rlabel metal3 s 0 76712 800 76832 6 ring0_trim_b[8]
port 561 nsew signal output
rlabel metal3 s 0 78752 800 78872 6 ring0_trim_b[9]
port 562 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 ring10_clk
port 563 nsew signal input
rlabel metal3 s 0 194624 800 194744 6 ring11_clk
port 564 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 ring12_clk
port 565 nsew signal input
rlabel metal3 s 99200 189184 100000 189304 6 ring13_clk
port 566 nsew signal input
rlabel metal3 s 99200 192312 100000 192432 6 ring14_clk
port 567 nsew signal input
rlabel metal3 s 0 196800 800 196920 6 ring15_clk
port 568 nsew signal input
rlabel metal3 s 99200 195304 100000 195424 6 ring16_clk
port 569 nsew signal input
rlabel metal2 s 98642 199200 98698 200000 6 ring17_clk
port 570 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 ring18_clk
port 571 nsew signal input
rlabel metal2 s 99470 199200 99526 200000 6 ring19_clk
port 572 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 ring1_clk
port 573 nsew signal input
rlabel metal3 s 0 181976 800 182096 6 ring1_clkmux[0]
port 574 nsew signal output
rlabel metal3 s 0 184152 800 184272 6 ring1_clkmux[1]
port 575 nsew signal output
rlabel metal3 s 0 186192 800 186312 6 ring1_clkmux[2]
port 576 nsew signal output
rlabel metal3 s 0 188368 800 188488 6 ring1_start
port 577 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 ring1_trim_a[0]
port 578 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 ring1_trim_a[10]
port 579 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 ring1_trim_a[11]
port 580 nsew signal output
rlabel metal3 s 0 152464 800 152584 6 ring1_trim_a[12]
port 581 nsew signal output
rlabel metal3 s 0 154640 800 154760 6 ring1_trim_a[13]
port 582 nsew signal output
rlabel metal3 s 0 156680 800 156800 6 ring1_trim_a[14]
port 583 nsew signal output
rlabel metal3 s 0 158856 800 158976 6 ring1_trim_a[15]
port 584 nsew signal output
rlabel metal3 s 0 160896 800 161016 6 ring1_trim_a[16]
port 585 nsew signal output
rlabel metal3 s 0 163072 800 163192 6 ring1_trim_a[17]
port 586 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 ring1_trim_a[18]
port 587 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 ring1_trim_a[19]
port 588 nsew signal output
rlabel metal3 s 0 129344 800 129464 6 ring1_trim_a[1]
port 589 nsew signal output
rlabel metal3 s 0 169328 800 169448 6 ring1_trim_a[20]
port 590 nsew signal output
rlabel metal3 s 0 171504 800 171624 6 ring1_trim_a[21]
port 591 nsew signal output
rlabel metal3 s 0 173544 800 173664 6 ring1_trim_a[22]
port 592 nsew signal output
rlabel metal3 s 0 175720 800 175840 6 ring1_trim_a[23]
port 593 nsew signal output
rlabel metal3 s 0 177760 800 177880 6 ring1_trim_a[24]
port 594 nsew signal output
rlabel metal3 s 0 179936 800 180056 6 ring1_trim_a[25]
port 595 nsew signal output
rlabel metal3 s 0 131520 800 131640 6 ring1_trim_a[2]
port 596 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 ring1_trim_a[3]
port 597 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 ring1_trim_a[4]
port 598 nsew signal output
rlabel metal3 s 0 137776 800 137896 6 ring1_trim_a[5]
port 599 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 ring1_trim_a[6]
port 600 nsew signal output
rlabel metal3 s 0 141992 800 142112 6 ring1_trim_a[7]
port 601 nsew signal output
rlabel metal3 s 0 144032 800 144152 6 ring1_trim_a[8]
port 602 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 ring1_trim_a[9]
port 603 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 ring20_clk
port 604 nsew signal input
rlabel metal3 s 0 198840 800 198960 6 ring21_clk
port 605 nsew signal input
rlabel metal3 s 99200 198432 100000 198552 6 ring22_clk
port 606 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 ring2_clk
port 607 nsew signal input
rlabel metal3 s 99200 173816 100000 173936 6 ring2_clkmux[0]
port 608 nsew signal output
rlabel metal3 s 99200 176808 100000 176928 6 ring2_clkmux[1]
port 609 nsew signal output
rlabel metal3 s 99200 179936 100000 180056 6 ring2_clkmux[2]
port 610 nsew signal output
rlabel metal3 s 99200 183064 100000 183184 6 ring2_start
port 611 nsew signal output
rlabel metal3 s 99200 1504 100000 1624 6 ring2_trim_a[0]
port 612 nsew signal output
rlabel metal3 s 99200 32240 100000 32360 6 ring2_trim_a[10]
port 613 nsew signal output
rlabel metal3 s 99200 35232 100000 35352 6 ring2_trim_a[11]
port 614 nsew signal output
rlabel metal3 s 99200 38360 100000 38480 6 ring2_trim_a[12]
port 615 nsew signal output
rlabel metal3 s 99200 41488 100000 41608 6 ring2_trim_a[13]
port 616 nsew signal output
rlabel metal3 s 99200 44480 100000 44600 6 ring2_trim_a[14]
port 617 nsew signal output
rlabel metal3 s 99200 47608 100000 47728 6 ring2_trim_a[15]
port 618 nsew signal output
rlabel metal3 s 99200 50736 100000 50856 6 ring2_trim_a[16]
port 619 nsew signal output
rlabel metal3 s 99200 53728 100000 53848 6 ring2_trim_a[17]
port 620 nsew signal output
rlabel metal3 s 99200 56856 100000 56976 6 ring2_trim_a[18]
port 621 nsew signal output
rlabel metal3 s 99200 59848 100000 59968 6 ring2_trim_a[19]
port 622 nsew signal output
rlabel metal3 s 99200 4496 100000 4616 6 ring2_trim_a[1]
port 623 nsew signal output
rlabel metal3 s 99200 62976 100000 63096 6 ring2_trim_a[20]
port 624 nsew signal output
rlabel metal3 s 99200 66104 100000 66224 6 ring2_trim_a[21]
port 625 nsew signal output
rlabel metal3 s 99200 69096 100000 69216 6 ring2_trim_a[22]
port 626 nsew signal output
rlabel metal3 s 99200 72224 100000 72344 6 ring2_trim_a[23]
port 627 nsew signal output
rlabel metal3 s 99200 75352 100000 75472 6 ring2_trim_a[24]
port 628 nsew signal output
rlabel metal3 s 99200 78344 100000 78464 6 ring2_trim_a[25]
port 629 nsew signal output
rlabel metal3 s 99200 81472 100000 81592 6 ring2_trim_a[26]
port 630 nsew signal output
rlabel metal3 s 99200 84600 100000 84720 6 ring2_trim_a[27]
port 631 nsew signal output
rlabel metal3 s 99200 7624 100000 7744 6 ring2_trim_a[2]
port 632 nsew signal output
rlabel metal3 s 99200 10616 100000 10736 6 ring2_trim_a[3]
port 633 nsew signal output
rlabel metal3 s 99200 13744 100000 13864 6 ring2_trim_a[4]
port 634 nsew signal output
rlabel metal3 s 99200 16872 100000 16992 6 ring2_trim_a[5]
port 635 nsew signal output
rlabel metal3 s 99200 19864 100000 19984 6 ring2_trim_a[6]
port 636 nsew signal output
rlabel metal3 s 99200 22992 100000 23112 6 ring2_trim_a[7]
port 637 nsew signal output
rlabel metal3 s 99200 26120 100000 26240 6 ring2_trim_a[8]
port 638 nsew signal output
rlabel metal3 s 99200 29112 100000 29232 6 ring2_trim_a[9]
port 639 nsew signal output
rlabel metal3 s 99200 87592 100000 87712 6 ring2_trim_b[0]
port 640 nsew signal output
rlabel metal3 s 99200 118328 100000 118448 6 ring2_trim_b[10]
port 641 nsew signal output
rlabel metal3 s 99200 121456 100000 121576 6 ring2_trim_b[11]
port 642 nsew signal output
rlabel metal3 s 99200 124584 100000 124704 6 ring2_trim_b[12]
port 643 nsew signal output
rlabel metal3 s 99200 127576 100000 127696 6 ring2_trim_b[13]
port 644 nsew signal output
rlabel metal3 s 99200 130704 100000 130824 6 ring2_trim_b[14]
port 645 nsew signal output
rlabel metal3 s 99200 133832 100000 133952 6 ring2_trim_b[15]
port 646 nsew signal output
rlabel metal3 s 99200 136824 100000 136944 6 ring2_trim_b[16]
port 647 nsew signal output
rlabel metal3 s 99200 139952 100000 140072 6 ring2_trim_b[17]
port 648 nsew signal output
rlabel metal3 s 99200 143080 100000 143200 6 ring2_trim_b[18]
port 649 nsew signal output
rlabel metal3 s 99200 146072 100000 146192 6 ring2_trim_b[19]
port 650 nsew signal output
rlabel metal3 s 99200 90720 100000 90840 6 ring2_trim_b[1]
port 651 nsew signal output
rlabel metal3 s 99200 149200 100000 149320 6 ring2_trim_b[20]
port 652 nsew signal output
rlabel metal3 s 99200 152192 100000 152312 6 ring2_trim_b[21]
port 653 nsew signal output
rlabel metal3 s 99200 155320 100000 155440 6 ring2_trim_b[22]
port 654 nsew signal output
rlabel metal3 s 99200 158448 100000 158568 6 ring2_trim_b[23]
port 655 nsew signal output
rlabel metal3 s 99200 161440 100000 161560 6 ring2_trim_b[24]
port 656 nsew signal output
rlabel metal3 s 99200 164568 100000 164688 6 ring2_trim_b[25]
port 657 nsew signal output
rlabel metal3 s 99200 167696 100000 167816 6 ring2_trim_b[26]
port 658 nsew signal output
rlabel metal3 s 99200 170688 100000 170808 6 ring2_trim_b[27]
port 659 nsew signal output
rlabel metal3 s 99200 93712 100000 93832 6 ring2_trim_b[2]
port 660 nsew signal output
rlabel metal3 s 99200 96840 100000 96960 6 ring2_trim_b[3]
port 661 nsew signal output
rlabel metal3 s 99200 99968 100000 100088 6 ring2_trim_b[4]
port 662 nsew signal output
rlabel metal3 s 99200 102960 100000 103080 6 ring2_trim_b[5]
port 663 nsew signal output
rlabel metal3 s 99200 106088 100000 106208 6 ring2_trim_b[6]
port 664 nsew signal output
rlabel metal3 s 99200 109216 100000 109336 6 ring2_trim_b[7]
port 665 nsew signal output
rlabel metal3 s 99200 112208 100000 112328 6 ring2_trim_b[8]
port 666 nsew signal output
rlabel metal3 s 99200 115336 100000 115456 6 ring2_trim_b[9]
port 667 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 ring3_clk
port 668 nsew signal input
rlabel metal2 s 96986 199200 97042 200000 6 ring4_clk
port 669 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 ring5_clk
port 670 nsew signal input
rlabel metal3 s 99200 186056 100000 186176 6 ring6_clk
port 671 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 ring7_clk
port 672 nsew signal input
rlabel metal3 s 0 192584 800 192704 6 ring8_clk
port 673 nsew signal input
rlabel metal2 s 97814 199200 97870 200000 6 ring9_clk
port 674 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 675 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 675 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 675 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 675 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 676 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 676 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 676 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 677 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 678 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 679 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wbs_adr_i[0]
port 680 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[10]
port 681 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[11]
port 682 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[12]
port 683 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[13]
port 684 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[14]
port 685 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[15]
port 686 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[16]
port 687 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[17]
port 688 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[18]
port 689 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[19]
port 690 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[1]
port 691 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[20]
port 692 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[21]
port 693 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[22]
port 694 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[23]
port 695 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[24]
port 696 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[25]
port 697 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[26]
port 698 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[27]
port 699 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[28]
port 700 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[29]
port 701 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 702 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[30]
port 703 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[31]
port 704 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[3]
port 705 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[4]
port 706 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[5]
port 707 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[6]
port 708 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_adr_i[7]
port 709 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[8]
port 710 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[9]
port 711 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 712 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 713 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[10]
port 714 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[11]
port 715 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[12]
port 716 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[13]
port 717 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[14]
port 718 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_i[15]
port 719 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[16]
port 720 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[17]
port 721 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[18]
port 722 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[19]
port 723 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_i[1]
port 724 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[20]
port 725 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[21]
port 726 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[22]
port 727 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[23]
port 728 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_i[24]
port 729 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[25]
port 730 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_i[26]
port 731 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[27]
port 732 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[28]
port 733 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_i[29]
port 734 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[2]
port 735 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[30]
port 736 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[31]
port 737 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 738 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[4]
port 739 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[5]
port 740 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[6]
port 741 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[7]
port 742 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[8]
port 743 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[9]
port 744 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 745 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[10]
port 746 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[11]
port 747 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[12]
port 748 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_o[13]
port 749 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[14]
port 750 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[15]
port 751 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[16]
port 752 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[17]
port 753 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[18]
port 754 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[19]
port 755 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[1]
port 756 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[20]
port 757 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_o[21]
port 758 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[22]
port 759 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[23]
port 760 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_o[24]
port 761 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[25]
port 762 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[26]
port 763 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[27]
port 764 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[28]
port 765 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[29]
port 766 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[2]
port 767 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_o[30]
port 768 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[31]
port 769 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_o[3]
port 770 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[4]
port 771 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_o[5]
port 772 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[6]
port 773 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[7]
port 774 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[8]
port 775 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[9]
port 776 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 777 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 778 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_sel_i[2]
port 779 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_sel_i[3]
port 780 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 781 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_we_i
port 782 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/digitalcore_macro/runs/digitalcore_macro/results/magic/digitalcore_macro.gds
string GDS_END 29455782
string GDS_START 770462
<< end >>

