magic
tech sky130A
magscale 1 2
timestamp 1641023160
<< obsli1 >>
rect 1104 2159 99147 197489
<< obsm1 >>
rect 106 1232 99898 197520
<< metal2 >>
rect 386 199200 442 200000
rect 1214 199200 1270 200000
rect 2042 199200 2098 200000
rect 2962 199200 3018 200000
rect 3790 199200 3846 200000
rect 4710 199200 4766 200000
rect 5538 199200 5594 200000
rect 6458 199200 6514 200000
rect 7286 199200 7342 200000
rect 8206 199200 8262 200000
rect 9034 199200 9090 200000
rect 9862 199200 9918 200000
rect 10782 199200 10838 200000
rect 11610 199200 11666 200000
rect 12530 199200 12586 200000
rect 13358 199200 13414 200000
rect 14278 199200 14334 200000
rect 15106 199200 15162 200000
rect 16026 199200 16082 200000
rect 16854 199200 16910 200000
rect 17774 199200 17830 200000
rect 18602 199200 18658 200000
rect 19430 199200 19486 200000
rect 20350 199200 20406 200000
rect 21178 199200 21234 200000
rect 22098 199200 22154 200000
rect 22926 199200 22982 200000
rect 23846 199200 23902 200000
rect 24674 199200 24730 200000
rect 25594 199200 25650 200000
rect 26422 199200 26478 200000
rect 27342 199200 27398 200000
rect 28170 199200 28226 200000
rect 28998 199200 29054 200000
rect 29918 199200 29974 200000
rect 30746 199200 30802 200000
rect 31666 199200 31722 200000
rect 32494 199200 32550 200000
rect 33414 199200 33470 200000
rect 34242 199200 34298 200000
rect 35162 199200 35218 200000
rect 35990 199200 36046 200000
rect 36818 199200 36874 200000
rect 37738 199200 37794 200000
rect 38566 199200 38622 200000
rect 39486 199200 39542 200000
rect 40314 199200 40370 200000
rect 41234 199200 41290 200000
rect 42062 199200 42118 200000
rect 42982 199200 43038 200000
rect 43810 199200 43866 200000
rect 44730 199200 44786 200000
rect 45558 199200 45614 200000
rect 46386 199200 46442 200000
rect 47306 199200 47362 200000
rect 48134 199200 48190 200000
rect 49054 199200 49110 200000
rect 49882 199200 49938 200000
rect 50802 199200 50858 200000
rect 51630 199200 51686 200000
rect 52550 199200 52606 200000
rect 53378 199200 53434 200000
rect 54298 199200 54354 200000
rect 55126 199200 55182 200000
rect 55954 199200 56010 200000
rect 56874 199200 56930 200000
rect 57702 199200 57758 200000
rect 58622 199200 58678 200000
rect 59450 199200 59506 200000
rect 60370 199200 60426 200000
rect 61198 199200 61254 200000
rect 62118 199200 62174 200000
rect 62946 199200 63002 200000
rect 63866 199200 63922 200000
rect 64694 199200 64750 200000
rect 65522 199200 65578 200000
rect 66442 199200 66498 200000
rect 67270 199200 67326 200000
rect 68190 199200 68246 200000
rect 69018 199200 69074 200000
rect 69938 199200 69994 200000
rect 70766 199200 70822 200000
rect 71686 199200 71742 200000
rect 72514 199200 72570 200000
rect 73342 199200 73398 200000
rect 74262 199200 74318 200000
rect 75090 199200 75146 200000
rect 76010 199200 76066 200000
rect 76838 199200 76894 200000
rect 77758 199200 77814 200000
rect 78586 199200 78642 200000
rect 79506 199200 79562 200000
rect 80334 199200 80390 200000
rect 81254 199200 81310 200000
rect 82082 199200 82138 200000
rect 82910 199200 82966 200000
rect 83830 199200 83886 200000
rect 84658 199200 84714 200000
rect 85578 199200 85634 200000
rect 86406 199200 86462 200000
rect 87326 199200 87382 200000
rect 88154 199200 88210 200000
rect 89074 199200 89130 200000
rect 89902 199200 89958 200000
rect 90822 199200 90878 200000
rect 91650 199200 91706 200000
rect 92478 199200 92534 200000
rect 93398 199200 93454 200000
rect 94226 199200 94282 200000
rect 95146 199200 95202 200000
rect 95974 199200 96030 200000
rect 96894 199200 96950 200000
rect 97722 199200 97778 200000
rect 98642 199200 98698 200000
rect 99470 199200 99526 200000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16026 0 16082 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18050 0 18106 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19890 0 19946 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51538 0 51594 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65522 0 65578 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 69938 0 69994 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 71962 0 72018 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75826 0 75882 800
rect 76010 0 76066 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77482 0 77538 800
rect 77666 0 77722 800
rect 77850 0 77906 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79506 0 79562 800
rect 79690 0 79746 800
rect 79874 0 79930 800
rect 80058 0 80114 800
rect 80242 0 80298 800
rect 80426 0 80482 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82082 0 82138 800
rect 82266 0 82322 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 83922 0 83978 800
rect 84106 0 84162 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86130 0 86186 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 87970 0 88026 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89810 0 89866 800
rect 89994 0 90050 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 94042 0 94098 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 199144 330 199200
rect 498 199144 1158 199200
rect 1326 199144 1986 199200
rect 2154 199144 2906 199200
rect 3074 199144 3734 199200
rect 3902 199144 4654 199200
rect 4822 199144 5482 199200
rect 5650 199144 6402 199200
rect 6570 199144 7230 199200
rect 7398 199144 8150 199200
rect 8318 199144 8978 199200
rect 9146 199144 9806 199200
rect 9974 199144 10726 199200
rect 10894 199144 11554 199200
rect 11722 199144 12474 199200
rect 12642 199144 13302 199200
rect 13470 199144 14222 199200
rect 14390 199144 15050 199200
rect 15218 199144 15970 199200
rect 16138 199144 16798 199200
rect 16966 199144 17718 199200
rect 17886 199144 18546 199200
rect 18714 199144 19374 199200
rect 19542 199144 20294 199200
rect 20462 199144 21122 199200
rect 21290 199144 22042 199200
rect 22210 199144 22870 199200
rect 23038 199144 23790 199200
rect 23958 199144 24618 199200
rect 24786 199144 25538 199200
rect 25706 199144 26366 199200
rect 26534 199144 27286 199200
rect 27454 199144 28114 199200
rect 28282 199144 28942 199200
rect 29110 199144 29862 199200
rect 30030 199144 30690 199200
rect 30858 199144 31610 199200
rect 31778 199144 32438 199200
rect 32606 199144 33358 199200
rect 33526 199144 34186 199200
rect 34354 199144 35106 199200
rect 35274 199144 35934 199200
rect 36102 199144 36762 199200
rect 36930 199144 37682 199200
rect 37850 199144 38510 199200
rect 38678 199144 39430 199200
rect 39598 199144 40258 199200
rect 40426 199144 41178 199200
rect 41346 199144 42006 199200
rect 42174 199144 42926 199200
rect 43094 199144 43754 199200
rect 43922 199144 44674 199200
rect 44842 199144 45502 199200
rect 45670 199144 46330 199200
rect 46498 199144 47250 199200
rect 47418 199144 48078 199200
rect 48246 199144 48998 199200
rect 49166 199144 49826 199200
rect 49994 199144 50746 199200
rect 50914 199144 51574 199200
rect 51742 199144 52494 199200
rect 52662 199144 53322 199200
rect 53490 199144 54242 199200
rect 54410 199144 55070 199200
rect 55238 199144 55898 199200
rect 56066 199144 56818 199200
rect 56986 199144 57646 199200
rect 57814 199144 58566 199200
rect 58734 199144 59394 199200
rect 59562 199144 60314 199200
rect 60482 199144 61142 199200
rect 61310 199144 62062 199200
rect 62230 199144 62890 199200
rect 63058 199144 63810 199200
rect 63978 199144 64638 199200
rect 64806 199144 65466 199200
rect 65634 199144 66386 199200
rect 66554 199144 67214 199200
rect 67382 199144 68134 199200
rect 68302 199144 68962 199200
rect 69130 199144 69882 199200
rect 70050 199144 70710 199200
rect 70878 199144 71630 199200
rect 71798 199144 72458 199200
rect 72626 199144 73286 199200
rect 73454 199144 74206 199200
rect 74374 199144 75034 199200
rect 75202 199144 75954 199200
rect 76122 199144 76782 199200
rect 76950 199144 77702 199200
rect 77870 199144 78530 199200
rect 78698 199144 79450 199200
rect 79618 199144 80278 199200
rect 80446 199144 81198 199200
rect 81366 199144 82026 199200
rect 82194 199144 82854 199200
rect 83022 199144 83774 199200
rect 83942 199144 84602 199200
rect 84770 199144 85522 199200
rect 85690 199144 86350 199200
rect 86518 199144 87270 199200
rect 87438 199144 88098 199200
rect 88266 199144 89018 199200
rect 89186 199144 89846 199200
rect 90014 199144 90766 199200
rect 90934 199144 91594 199200
rect 91762 199144 92422 199200
rect 92590 199144 93342 199200
rect 93510 199144 94170 199200
rect 94338 199144 95090 199200
rect 95258 199144 95918 199200
rect 96086 199144 96838 199200
rect 97006 199144 97666 199200
rect 97834 199144 98586 199200
rect 98754 199144 99414 199200
rect 99582 199144 99892 199200
rect 112 856 99892 199144
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 974 856
rect 1142 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 1986 856
rect 2154 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 2998 856
rect 3166 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4010 856
rect 4178 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4838 856
rect 5006 800 5022 856
rect 5190 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5850 856
rect 6018 800 6034 856
rect 6202 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7046 856
rect 7214 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7874 856
rect 8042 800 8058 856
rect 8226 800 8334 856
rect 8502 800 8518 856
rect 8686 800 8702 856
rect 8870 800 8886 856
rect 9054 800 9070 856
rect 9238 800 9346 856
rect 9514 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10082 856
rect 10250 800 10266 856
rect 10434 800 10542 856
rect 10710 800 10726 856
rect 10894 800 10910 856
rect 11078 800 11094 856
rect 11262 800 11278 856
rect 11446 800 11554 856
rect 11722 800 11738 856
rect 11906 800 11922 856
rect 12090 800 12106 856
rect 12274 800 12290 856
rect 12458 800 12566 856
rect 12734 800 12750 856
rect 12918 800 12934 856
rect 13102 800 13118 856
rect 13286 800 13302 856
rect 13470 800 13578 856
rect 13746 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14130 856
rect 14298 800 14314 856
rect 14482 800 14590 856
rect 14758 800 14774 856
rect 14942 800 14958 856
rect 15126 800 15142 856
rect 15310 800 15326 856
rect 15494 800 15602 856
rect 15770 800 15786 856
rect 15954 800 15970 856
rect 16138 800 16154 856
rect 16322 800 16338 856
rect 16506 800 16614 856
rect 16782 800 16798 856
rect 16966 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17350 856
rect 17518 800 17626 856
rect 17794 800 17810 856
rect 17978 800 17994 856
rect 18162 800 18178 856
rect 18346 800 18362 856
rect 18530 800 18638 856
rect 18806 800 18822 856
rect 18990 800 19006 856
rect 19174 800 19190 856
rect 19358 800 19374 856
rect 19542 800 19650 856
rect 19818 800 19834 856
rect 20002 800 20018 856
rect 20186 800 20202 856
rect 20370 800 20386 856
rect 20554 800 20570 856
rect 20738 800 20846 856
rect 21014 800 21030 856
rect 21198 800 21214 856
rect 21382 800 21398 856
rect 21566 800 21582 856
rect 21750 800 21858 856
rect 22026 800 22042 856
rect 22210 800 22226 856
rect 22394 800 22410 856
rect 22578 800 22594 856
rect 22762 800 22870 856
rect 23038 800 23054 856
rect 23222 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24250 856
rect 24418 800 24434 856
rect 24602 800 24618 856
rect 24786 800 24894 856
rect 25062 800 25078 856
rect 25246 800 25262 856
rect 25430 800 25446 856
rect 25614 800 25630 856
rect 25798 800 25906 856
rect 26074 800 26090 856
rect 26258 800 26274 856
rect 26442 800 26458 856
rect 26626 800 26642 856
rect 26810 800 26918 856
rect 27086 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27654 856
rect 27822 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28298 856
rect 28466 800 28482 856
rect 28650 800 28666 856
rect 28834 800 28942 856
rect 29110 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29494 856
rect 29662 800 29678 856
rect 29846 800 29954 856
rect 30122 800 30138 856
rect 30306 800 30322 856
rect 30490 800 30506 856
rect 30674 800 30690 856
rect 30858 800 30874 856
rect 31042 800 31150 856
rect 31318 800 31334 856
rect 31502 800 31518 856
rect 31686 800 31702 856
rect 31870 800 31886 856
rect 32054 800 32162 856
rect 32330 800 32346 856
rect 32514 800 32530 856
rect 32698 800 32714 856
rect 32882 800 32898 856
rect 33066 800 33174 856
rect 33342 800 33358 856
rect 33526 800 33542 856
rect 33710 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34554 856
rect 34722 800 34738 856
rect 34906 800 34922 856
rect 35090 800 35198 856
rect 35366 800 35382 856
rect 35550 800 35566 856
rect 35734 800 35750 856
rect 35918 800 35934 856
rect 36102 800 36210 856
rect 36378 800 36394 856
rect 36562 800 36578 856
rect 36746 800 36762 856
rect 36930 800 36946 856
rect 37114 800 37222 856
rect 37390 800 37406 856
rect 37574 800 37590 856
rect 37758 800 37774 856
rect 37942 800 37958 856
rect 38126 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38602 856
rect 38770 800 38786 856
rect 38954 800 38970 856
rect 39138 800 39246 856
rect 39414 800 39430 856
rect 39598 800 39614 856
rect 39782 800 39798 856
rect 39966 800 39982 856
rect 40150 800 40166 856
rect 40334 800 40442 856
rect 40610 800 40626 856
rect 40794 800 40810 856
rect 40978 800 40994 856
rect 41162 800 41178 856
rect 41346 800 41454 856
rect 41622 800 41638 856
rect 41806 800 41822 856
rect 41990 800 42006 856
rect 42174 800 42190 856
rect 42358 800 42466 856
rect 42634 800 42650 856
rect 42818 800 42834 856
rect 43002 800 43018 856
rect 43186 800 43202 856
rect 43370 800 43478 856
rect 43646 800 43662 856
rect 43830 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44674 856
rect 44842 800 44858 856
rect 45026 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45502 856
rect 45670 800 45686 856
rect 45854 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46238 856
rect 46406 800 46514 856
rect 46682 800 46698 856
rect 46866 800 46882 856
rect 47050 800 47066 856
rect 47234 800 47250 856
rect 47418 800 47526 856
rect 47694 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48262 856
rect 48430 800 48538 856
rect 48706 800 48722 856
rect 48890 800 48906 856
rect 49074 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49550 856
rect 49718 800 49734 856
rect 49902 800 49918 856
rect 50086 800 50102 856
rect 50270 800 50286 856
rect 50454 800 50470 856
rect 50638 800 50746 856
rect 50914 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51298 856
rect 51466 800 51482 856
rect 51650 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52126 856
rect 52294 800 52310 856
rect 52478 800 52494 856
rect 52662 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53138 856
rect 53306 800 53322 856
rect 53490 800 53506 856
rect 53674 800 53782 856
rect 53950 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54334 856
rect 54502 800 54518 856
rect 54686 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55162 856
rect 55330 800 55346 856
rect 55514 800 55530 856
rect 55698 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56174 856
rect 56342 800 56358 856
rect 56526 800 56542 856
rect 56710 800 56818 856
rect 56986 800 57002 856
rect 57170 800 57186 856
rect 57354 800 57370 856
rect 57538 800 57554 856
rect 57722 800 57830 856
rect 57998 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58382 856
rect 58550 800 58566 856
rect 58734 800 58842 856
rect 59010 800 59026 856
rect 59194 800 59210 856
rect 59378 800 59394 856
rect 59562 800 59578 856
rect 59746 800 59854 856
rect 60022 800 60038 856
rect 60206 800 60222 856
rect 60390 800 60406 856
rect 60574 800 60590 856
rect 60758 800 60774 856
rect 60942 800 61050 856
rect 61218 800 61234 856
rect 61402 800 61418 856
rect 61586 800 61602 856
rect 61770 800 61786 856
rect 61954 800 62062 856
rect 62230 800 62246 856
rect 62414 800 62430 856
rect 62598 800 62614 856
rect 62782 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63258 856
rect 63426 800 63442 856
rect 63610 800 63626 856
rect 63794 800 63810 856
rect 63978 800 64086 856
rect 64254 800 64270 856
rect 64438 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64822 856
rect 64990 800 65098 856
rect 65266 800 65282 856
rect 65450 800 65466 856
rect 65634 800 65650 856
rect 65818 800 65834 856
rect 66002 800 66110 856
rect 66278 800 66294 856
rect 66462 800 66478 856
rect 66646 800 66662 856
rect 66830 800 66846 856
rect 67014 800 67122 856
rect 67290 800 67306 856
rect 67474 800 67490 856
rect 67658 800 67674 856
rect 67842 800 67858 856
rect 68026 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68686 856
rect 68854 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69330 856
rect 69498 800 69514 856
rect 69682 800 69698 856
rect 69866 800 69882 856
rect 70050 800 70066 856
rect 70234 800 70342 856
rect 70510 800 70526 856
rect 70694 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71078 856
rect 71246 800 71354 856
rect 71522 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71906 856
rect 72074 800 72090 856
rect 72258 800 72366 856
rect 72534 800 72550 856
rect 72718 800 72734 856
rect 72902 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73378 856
rect 73546 800 73562 856
rect 73730 800 73746 856
rect 73914 800 73930 856
rect 74098 800 74114 856
rect 74282 800 74390 856
rect 74558 800 74574 856
rect 74742 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75126 856
rect 75294 800 75402 856
rect 75570 800 75586 856
rect 75754 800 75770 856
rect 75938 800 75954 856
rect 76122 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76598 856
rect 76766 800 76782 856
rect 76950 800 76966 856
rect 77134 800 77150 856
rect 77318 800 77426 856
rect 77594 800 77610 856
rect 77778 800 77794 856
rect 77962 800 77978 856
rect 78146 800 78162 856
rect 78330 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78806 856
rect 78974 800 78990 856
rect 79158 800 79174 856
rect 79342 800 79450 856
rect 79618 800 79634 856
rect 79802 800 79818 856
rect 79986 800 80002 856
rect 80170 800 80186 856
rect 80354 800 80370 856
rect 80538 800 80646 856
rect 80814 800 80830 856
rect 80998 800 81014 856
rect 81182 800 81198 856
rect 81366 800 81382 856
rect 81550 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82026 856
rect 82194 800 82210 856
rect 82378 800 82394 856
rect 82562 800 82670 856
rect 82838 800 82854 856
rect 83022 800 83038 856
rect 83206 800 83222 856
rect 83390 800 83406 856
rect 83574 800 83682 856
rect 83850 800 83866 856
rect 84034 800 84050 856
rect 84218 800 84234 856
rect 84402 800 84418 856
rect 84586 800 84694 856
rect 84862 800 84878 856
rect 85046 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85430 856
rect 85598 800 85706 856
rect 85874 800 85890 856
rect 86058 800 86074 856
rect 86242 800 86258 856
rect 86426 800 86442 856
rect 86610 800 86718 856
rect 86886 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87730 856
rect 87898 800 87914 856
rect 88082 800 88098 856
rect 88266 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89110 856
rect 89278 800 89294 856
rect 89462 800 89478 856
rect 89646 800 89754 856
rect 89922 800 89938 856
rect 90106 800 90122 856
rect 90290 800 90306 856
rect 90474 800 90490 856
rect 90658 800 90674 856
rect 90842 800 90950 856
rect 91118 800 91134 856
rect 91302 800 91318 856
rect 91486 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91962 856
rect 92130 800 92146 856
rect 92314 800 92330 856
rect 92498 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92974 856
rect 93142 800 93158 856
rect 93326 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93710 856
rect 93878 800 93986 856
rect 94154 800 94170 856
rect 94338 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94998 856
rect 95166 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 96010 856
rect 96178 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 98034 856
rect 98202 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 99046 856
rect 99214 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 198840 800 198960
rect 99200 198432 100000 198552
rect 0 196664 800 196784
rect 99200 195304 100000 195424
rect 0 194488 800 194608
rect 0 192312 800 192432
rect 99200 192176 100000 192296
rect 0 190136 800 190256
rect 99200 189048 100000 189168
rect 0 188096 800 188216
rect 0 185920 800 186040
rect 99200 185920 100000 186040
rect 0 183744 800 183864
rect 99200 182792 100000 182912
rect 0 181568 800 181688
rect 99200 179664 100000 179784
rect 0 179392 800 179512
rect 0 177352 800 177472
rect 99200 176536 100000 176656
rect 0 175176 800 175296
rect 99200 173408 100000 173528
rect 0 173000 800 173120
rect 0 170824 800 170944
rect 99200 170280 100000 170400
rect 0 168648 800 168768
rect 99200 167152 100000 167272
rect 0 166472 800 166592
rect 0 164432 800 164552
rect 99200 164024 100000 164144
rect 0 162256 800 162376
rect 99200 160896 100000 161016
rect 0 160080 800 160200
rect 0 157904 800 158024
rect 99200 157768 100000 157888
rect 0 155728 800 155848
rect 99200 154640 100000 154760
rect 0 153688 800 153808
rect 0 151512 800 151632
rect 99200 151512 100000 151632
rect 0 149336 800 149456
rect 99200 148384 100000 148504
rect 0 147160 800 147280
rect 99200 145256 100000 145376
rect 0 144984 800 145104
rect 0 142808 800 142928
rect 99200 142128 100000 142248
rect 0 140768 800 140888
rect 99200 139000 100000 139120
rect 0 138592 800 138712
rect 0 136416 800 136536
rect 99200 135872 100000 135992
rect 0 134240 800 134360
rect 99200 132744 100000 132864
rect 0 132064 800 132184
rect 0 130024 800 130144
rect 99200 129616 100000 129736
rect 0 127848 800 127968
rect 99200 126488 100000 126608
rect 0 125672 800 125792
rect 0 123496 800 123616
rect 99200 123360 100000 123480
rect 0 121320 800 121440
rect 99200 120232 100000 120352
rect 0 119144 800 119264
rect 0 117104 800 117224
rect 99200 117104 100000 117224
rect 0 114928 800 115048
rect 99200 113976 100000 114096
rect 0 112752 800 112872
rect 99200 110848 100000 110968
rect 0 110576 800 110696
rect 0 108400 800 108520
rect 99200 107720 100000 107840
rect 0 106360 800 106480
rect 99200 104592 100000 104712
rect 0 104184 800 104304
rect 0 102008 800 102128
rect 99200 101464 100000 101584
rect 0 99832 800 99952
rect 99200 98336 100000 98456
rect 0 97656 800 97776
rect 0 95480 800 95600
rect 99200 95208 100000 95328
rect 0 93440 800 93560
rect 99200 92080 100000 92200
rect 0 91264 800 91384
rect 0 89088 800 89208
rect 99200 88952 100000 89072
rect 0 86912 800 87032
rect 99200 85824 100000 85944
rect 0 84736 800 84856
rect 0 82696 800 82816
rect 99200 82696 100000 82816
rect 0 80520 800 80640
rect 99200 79568 100000 79688
rect 0 78344 800 78464
rect 99200 76440 100000 76560
rect 0 76168 800 76288
rect 0 73992 800 74112
rect 99200 73312 100000 73432
rect 0 71816 800 71936
rect 99200 70184 100000 70304
rect 0 69776 800 69896
rect 0 67600 800 67720
rect 99200 67056 100000 67176
rect 0 65424 800 65544
rect 99200 63928 100000 64048
rect 0 63248 800 63368
rect 0 61072 800 61192
rect 99200 60800 100000 60920
rect 0 59032 800 59152
rect 99200 57672 100000 57792
rect 0 56856 800 56976
rect 0 54680 800 54800
rect 99200 54544 100000 54664
rect 0 52504 800 52624
rect 99200 51416 100000 51536
rect 0 50328 800 50448
rect 0 48152 800 48272
rect 99200 48288 100000 48408
rect 0 46112 800 46232
rect 99200 45160 100000 45280
rect 0 43936 800 44056
rect 99200 42032 100000 42152
rect 0 41760 800 41880
rect 0 39584 800 39704
rect 99200 38904 100000 39024
rect 0 37408 800 37528
rect 99200 35776 100000 35896
rect 0 35368 800 35488
rect 0 33192 800 33312
rect 99200 32648 100000 32768
rect 0 31016 800 31136
rect 99200 29520 100000 29640
rect 0 28840 800 28960
rect 0 26664 800 26784
rect 99200 26392 100000 26512
rect 0 24488 800 24608
rect 99200 23264 100000 23384
rect 0 22448 800 22568
rect 0 20272 800 20392
rect 99200 20136 100000 20256
rect 0 18096 800 18216
rect 99200 17008 100000 17128
rect 0 15920 800 16040
rect 0 13744 800 13864
rect 99200 13880 100000 14000
rect 0 11704 800 11824
rect 99200 10752 100000 10872
rect 0 9528 800 9648
rect 99200 7624 100000 7744
rect 0 7352 800 7472
rect 0 5176 800 5296
rect 99200 4496 100000 4616
rect 0 3000 800 3120
rect 99200 1504 100000 1624
rect 0 960 800 1080
<< obsm3 >>
rect 880 198760 99200 198933
rect 800 198632 99200 198760
rect 800 198352 99120 198632
rect 800 196864 99200 198352
rect 880 196584 99200 196864
rect 800 195504 99200 196584
rect 800 195224 99120 195504
rect 800 194688 99200 195224
rect 880 194408 99200 194688
rect 800 192512 99200 194408
rect 880 192376 99200 192512
rect 880 192232 99120 192376
rect 800 192096 99120 192232
rect 800 190336 99200 192096
rect 880 190056 99200 190336
rect 800 189248 99200 190056
rect 800 188968 99120 189248
rect 800 188296 99200 188968
rect 880 188016 99200 188296
rect 800 186120 99200 188016
rect 880 185840 99120 186120
rect 800 183944 99200 185840
rect 880 183664 99200 183944
rect 800 182992 99200 183664
rect 800 182712 99120 182992
rect 800 181768 99200 182712
rect 880 181488 99200 181768
rect 800 179864 99200 181488
rect 800 179592 99120 179864
rect 880 179584 99120 179592
rect 880 179312 99200 179584
rect 800 177552 99200 179312
rect 880 177272 99200 177552
rect 800 176736 99200 177272
rect 800 176456 99120 176736
rect 800 175376 99200 176456
rect 880 175096 99200 175376
rect 800 173608 99200 175096
rect 800 173328 99120 173608
rect 800 173200 99200 173328
rect 880 172920 99200 173200
rect 800 171024 99200 172920
rect 880 170744 99200 171024
rect 800 170480 99200 170744
rect 800 170200 99120 170480
rect 800 168848 99200 170200
rect 880 168568 99200 168848
rect 800 167352 99200 168568
rect 800 167072 99120 167352
rect 800 166672 99200 167072
rect 880 166392 99200 166672
rect 800 164632 99200 166392
rect 880 164352 99200 164632
rect 800 164224 99200 164352
rect 800 163944 99120 164224
rect 800 162456 99200 163944
rect 880 162176 99200 162456
rect 800 161096 99200 162176
rect 800 160816 99120 161096
rect 800 160280 99200 160816
rect 880 160000 99200 160280
rect 800 158104 99200 160000
rect 880 157968 99200 158104
rect 880 157824 99120 157968
rect 800 157688 99120 157824
rect 800 155928 99200 157688
rect 880 155648 99200 155928
rect 800 154840 99200 155648
rect 800 154560 99120 154840
rect 800 153888 99200 154560
rect 880 153608 99200 153888
rect 800 151712 99200 153608
rect 880 151432 99120 151712
rect 800 149536 99200 151432
rect 880 149256 99200 149536
rect 800 148584 99200 149256
rect 800 148304 99120 148584
rect 800 147360 99200 148304
rect 880 147080 99200 147360
rect 800 145456 99200 147080
rect 800 145184 99120 145456
rect 880 145176 99120 145184
rect 880 144904 99200 145176
rect 800 143008 99200 144904
rect 880 142728 99200 143008
rect 800 142328 99200 142728
rect 800 142048 99120 142328
rect 800 140968 99200 142048
rect 880 140688 99200 140968
rect 800 139200 99200 140688
rect 800 138920 99120 139200
rect 800 138792 99200 138920
rect 880 138512 99200 138792
rect 800 136616 99200 138512
rect 880 136336 99200 136616
rect 800 136072 99200 136336
rect 800 135792 99120 136072
rect 800 134440 99200 135792
rect 880 134160 99200 134440
rect 800 132944 99200 134160
rect 800 132664 99120 132944
rect 800 132264 99200 132664
rect 880 131984 99200 132264
rect 800 130224 99200 131984
rect 880 129944 99200 130224
rect 800 129816 99200 129944
rect 800 129536 99120 129816
rect 800 128048 99200 129536
rect 880 127768 99200 128048
rect 800 126688 99200 127768
rect 800 126408 99120 126688
rect 800 125872 99200 126408
rect 880 125592 99200 125872
rect 800 123696 99200 125592
rect 880 123560 99200 123696
rect 880 123416 99120 123560
rect 800 123280 99120 123416
rect 800 121520 99200 123280
rect 880 121240 99200 121520
rect 800 120432 99200 121240
rect 800 120152 99120 120432
rect 800 119344 99200 120152
rect 880 119064 99200 119344
rect 800 117304 99200 119064
rect 880 117024 99120 117304
rect 800 115128 99200 117024
rect 880 114848 99200 115128
rect 800 114176 99200 114848
rect 800 113896 99120 114176
rect 800 112952 99200 113896
rect 880 112672 99200 112952
rect 800 111048 99200 112672
rect 800 110776 99120 111048
rect 880 110768 99120 110776
rect 880 110496 99200 110768
rect 800 108600 99200 110496
rect 880 108320 99200 108600
rect 800 107920 99200 108320
rect 800 107640 99120 107920
rect 800 106560 99200 107640
rect 880 106280 99200 106560
rect 800 104792 99200 106280
rect 800 104512 99120 104792
rect 800 104384 99200 104512
rect 880 104104 99200 104384
rect 800 102208 99200 104104
rect 880 101928 99200 102208
rect 800 101664 99200 101928
rect 800 101384 99120 101664
rect 800 100032 99200 101384
rect 880 99752 99200 100032
rect 800 98536 99200 99752
rect 800 98256 99120 98536
rect 800 97856 99200 98256
rect 880 97576 99200 97856
rect 800 95680 99200 97576
rect 880 95408 99200 95680
rect 880 95400 99120 95408
rect 800 95128 99120 95400
rect 800 93640 99200 95128
rect 880 93360 99200 93640
rect 800 92280 99200 93360
rect 800 92000 99120 92280
rect 800 91464 99200 92000
rect 880 91184 99200 91464
rect 800 89288 99200 91184
rect 880 89152 99200 89288
rect 880 89008 99120 89152
rect 800 88872 99120 89008
rect 800 87112 99200 88872
rect 880 86832 99200 87112
rect 800 86024 99200 86832
rect 800 85744 99120 86024
rect 800 84936 99200 85744
rect 880 84656 99200 84936
rect 800 82896 99200 84656
rect 880 82616 99120 82896
rect 800 80720 99200 82616
rect 880 80440 99200 80720
rect 800 79768 99200 80440
rect 800 79488 99120 79768
rect 800 78544 99200 79488
rect 880 78264 99200 78544
rect 800 76640 99200 78264
rect 800 76368 99120 76640
rect 880 76360 99120 76368
rect 880 76088 99200 76360
rect 800 74192 99200 76088
rect 880 73912 99200 74192
rect 800 73512 99200 73912
rect 800 73232 99120 73512
rect 800 72016 99200 73232
rect 880 71736 99200 72016
rect 800 70384 99200 71736
rect 800 70104 99120 70384
rect 800 69976 99200 70104
rect 880 69696 99200 69976
rect 800 67800 99200 69696
rect 880 67520 99200 67800
rect 800 67256 99200 67520
rect 800 66976 99120 67256
rect 800 65624 99200 66976
rect 880 65344 99200 65624
rect 800 64128 99200 65344
rect 800 63848 99120 64128
rect 800 63448 99200 63848
rect 880 63168 99200 63448
rect 800 61272 99200 63168
rect 880 61000 99200 61272
rect 880 60992 99120 61000
rect 800 60720 99120 60992
rect 800 59232 99200 60720
rect 880 58952 99200 59232
rect 800 57872 99200 58952
rect 800 57592 99120 57872
rect 800 57056 99200 57592
rect 880 56776 99200 57056
rect 800 54880 99200 56776
rect 880 54744 99200 54880
rect 880 54600 99120 54744
rect 800 54464 99120 54600
rect 800 52704 99200 54464
rect 880 52424 99200 52704
rect 800 51616 99200 52424
rect 800 51336 99120 51616
rect 800 50528 99200 51336
rect 880 50248 99200 50528
rect 800 48488 99200 50248
rect 800 48352 99120 48488
rect 880 48208 99120 48352
rect 880 48072 99200 48208
rect 800 46312 99200 48072
rect 880 46032 99200 46312
rect 800 45360 99200 46032
rect 800 45080 99120 45360
rect 800 44136 99200 45080
rect 880 43856 99200 44136
rect 800 42232 99200 43856
rect 800 41960 99120 42232
rect 880 41952 99120 41960
rect 880 41680 99200 41952
rect 800 39784 99200 41680
rect 880 39504 99200 39784
rect 800 39104 99200 39504
rect 800 38824 99120 39104
rect 800 37608 99200 38824
rect 880 37328 99200 37608
rect 800 35976 99200 37328
rect 800 35696 99120 35976
rect 800 35568 99200 35696
rect 880 35288 99200 35568
rect 800 33392 99200 35288
rect 880 33112 99200 33392
rect 800 32848 99200 33112
rect 800 32568 99120 32848
rect 800 31216 99200 32568
rect 880 30936 99200 31216
rect 800 29720 99200 30936
rect 800 29440 99120 29720
rect 800 29040 99200 29440
rect 880 28760 99200 29040
rect 800 26864 99200 28760
rect 880 26592 99200 26864
rect 880 26584 99120 26592
rect 800 26312 99120 26584
rect 800 24688 99200 26312
rect 880 24408 99200 24688
rect 800 23464 99200 24408
rect 800 23184 99120 23464
rect 800 22648 99200 23184
rect 880 22368 99200 22648
rect 800 20472 99200 22368
rect 880 20336 99200 20472
rect 880 20192 99120 20336
rect 800 20056 99120 20192
rect 800 18296 99200 20056
rect 880 18016 99200 18296
rect 800 17208 99200 18016
rect 800 16928 99120 17208
rect 800 16120 99200 16928
rect 880 15840 99200 16120
rect 800 14080 99200 15840
rect 800 13944 99120 14080
rect 880 13800 99120 13944
rect 880 13664 99200 13800
rect 800 11904 99200 13664
rect 880 11624 99200 11904
rect 800 10952 99200 11624
rect 800 10672 99120 10952
rect 800 9728 99200 10672
rect 880 9448 99200 9728
rect 800 7824 99200 9448
rect 800 7552 99120 7824
rect 880 7544 99120 7552
rect 880 7272 99200 7544
rect 800 5376 99200 7272
rect 880 5096 99200 5376
rect 800 4696 99200 5096
rect 800 4416 99120 4696
rect 800 3200 99200 4416
rect 880 2920 99200 3200
rect 800 1704 99200 2920
rect 800 1424 99120 1704
rect 800 1160 99200 1424
rect 880 987 99200 1160
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
<< obsm4 >>
rect 1715 2483 4128 192677
rect 4608 2483 19488 192677
rect 19968 2483 34848 192677
rect 35328 2483 43917 192677
<< labels >>
rlabel metal2 s 386 199200 442 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26422 199200 26478 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 28998 199200 29054 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31666 199200 31722 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34242 199200 34298 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 36818 199200 36874 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39486 199200 39542 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42062 199200 42118 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 44730 199200 44786 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47306 199200 47362 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 49882 199200 49938 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 199200 3018 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 52550 199200 52606 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55126 199200 55182 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57702 199200 57758 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60370 199200 60426 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 62946 199200 63002 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 65522 199200 65578 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68190 199200 68246 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70766 199200 70822 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73342 199200 73398 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76010 199200 76066 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5538 199200 5594 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 78586 199200 78642 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81254 199200 81310 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 83830 199200 83886 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 86406 199200 86462 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89074 199200 89130 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 91650 199200 91706 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 94226 199200 94282 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 96894 199200 96950 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 199200 8262 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10782 199200 10838 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13358 199200 13414 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16026 199200 16082 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18602 199200 18658 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21178 199200 21234 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23846 199200 23902 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 199200 1270 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27342 199200 27398 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 29918 199200 29974 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32494 199200 32550 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35162 199200 35218 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 37738 199200 37794 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40314 199200 40370 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 42982 199200 43038 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45558 199200 45614 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48134 199200 48190 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 50802 199200 50858 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3790 199200 3846 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53378 199200 53434 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 55954 199200 56010 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 58622 199200 58678 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61198 199200 61254 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 63866 199200 63922 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66442 199200 66498 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69018 199200 69074 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 71686 199200 71742 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74262 199200 74318 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 76838 199200 76894 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 199200 6514 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 79506 199200 79562 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82082 199200 82138 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 84658 199200 84714 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 87326 199200 87382 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 89902 199200 89958 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 92478 199200 92534 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95146 199200 95202 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 97722 199200 97778 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9034 199200 9090 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11610 199200 11666 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14278 199200 14334 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 16854 199200 16910 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19430 199200 19486 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22098 199200 22154 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24674 199200 24730 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2042 199200 2098 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28170 199200 28226 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 30746 199200 30802 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33414 199200 33470 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 35990 199200 36046 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38566 199200 38622 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41234 199200 41290 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 43810 199200 43866 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46386 199200 46442 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49054 199200 49110 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 51630 199200 51686 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 199200 4766 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54298 199200 54354 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 56874 199200 56930 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 59450 199200 59506 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62118 199200 62174 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 64694 199200 64750 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67270 199200 67326 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 69938 199200 69994 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 72514 199200 72570 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75090 199200 75146 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 77758 199200 77814 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7286 199200 7342 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 80334 199200 80390 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 82910 199200 82966 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 85578 199200 85634 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88154 199200 88210 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 90822 199200 90878 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 93398 199200 93454 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 95974 199200 96030 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 98642 199200 98698 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9862 199200 9918 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12530 199200 12586 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15106 199200 15162 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17774 199200 17830 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20350 199200 20406 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22926 199200 22982 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25594 199200 25650 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 0 194488 800 194608 6 ring0_clk
port 502 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 ring0_clkmux[0]
port 503 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 ring0_clkmux[1]
port 504 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 ring0_clkmux[2]
port 505 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 ring0_start
port 506 nsew signal output
rlabel metal3 s 0 960 800 1080 6 ring0_trim_a[0]
port 507 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 ring0_trim_a[10]
port 508 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 ring0_trim_a[11]
port 509 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 ring0_trim_a[12]
port 510 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 ring0_trim_a[13]
port 511 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 ring0_trim_a[14]
port 512 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 ring0_trim_a[15]
port 513 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 ring0_trim_a[16]
port 514 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 ring0_trim_a[17]
port 515 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 ring0_trim_a[18]
port 516 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 ring0_trim_a[19]
port 517 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 ring0_trim_a[1]
port 518 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 ring0_trim_a[20]
port 519 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 ring0_trim_a[21]
port 520 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 ring0_trim_a[22]
port 521 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 ring0_trim_a[23]
port 522 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 ring0_trim_a[24]
port 523 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 ring0_trim_a[25]
port 524 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 ring0_trim_a[26]
port 525 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 ring0_trim_a[27]
port 526 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 ring0_trim_a[2]
port 527 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 ring0_trim_a[3]
port 528 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 ring0_trim_a[4]
port 529 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 ring0_trim_a[5]
port 530 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 ring0_trim_a[6]
port 531 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 ring0_trim_a[7]
port 532 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 ring0_trim_a[8]
port 533 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 ring0_trim_a[9]
port 534 nsew signal output
rlabel metal3 s 0 61072 800 61192 6 ring0_trim_b[0]
port 535 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 ring0_trim_b[10]
port 536 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 ring0_trim_b[11]
port 537 nsew signal output
rlabel metal3 s 0 86912 800 87032 6 ring0_trim_b[12]
port 538 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 ring0_trim_b[13]
port 539 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 ring0_trim_b[14]
port 540 nsew signal output
rlabel metal3 s 0 93440 800 93560 6 ring0_trim_b[15]
port 541 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 ring0_trim_b[16]
port 542 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 ring0_trim_b[17]
port 543 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 ring0_trim_b[18]
port 544 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 ring0_trim_b[19]
port 545 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 ring0_trim_b[1]
port 546 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 ring0_trim_b[20]
port 547 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 ring0_trim_b[21]
port 548 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 ring0_trim_b[22]
port 549 nsew signal output
rlabel metal3 s 0 110576 800 110696 6 ring0_trim_b[23]
port 550 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 ring0_trim_b[24]
port 551 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 ring0_trim_b[25]
port 552 nsew signal output
rlabel metal3 s 0 117104 800 117224 6 ring0_trim_b[26]
port 553 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 ring0_trim_b[27]
port 554 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 ring0_trim_b[2]
port 555 nsew signal output
rlabel metal3 s 0 67600 800 67720 6 ring0_trim_b[3]
port 556 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 ring0_trim_b[4]
port 557 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 ring0_trim_b[5]
port 558 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 ring0_trim_b[6]
port 559 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 ring0_trim_b[7]
port 560 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 ring0_trim_b[8]
port 561 nsew signal output
rlabel metal3 s 0 80520 800 80640 6 ring0_trim_b[9]
port 562 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 ring1_clk
port 563 nsew signal input
rlabel metal3 s 0 185920 800 186040 6 ring1_clkmux[0]
port 564 nsew signal output
rlabel metal3 s 0 188096 800 188216 6 ring1_clkmux[1]
port 565 nsew signal output
rlabel metal3 s 0 190136 800 190256 6 ring1_clkmux[2]
port 566 nsew signal output
rlabel metal3 s 0 192312 800 192432 6 ring1_start
port 567 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 ring1_trim_a[0]
port 568 nsew signal output
rlabel metal3 s 0 151512 800 151632 6 ring1_trim_a[10]
port 569 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 ring1_trim_a[11]
port 570 nsew signal output
rlabel metal3 s 0 155728 800 155848 6 ring1_trim_a[12]
port 571 nsew signal output
rlabel metal3 s 0 157904 800 158024 6 ring1_trim_a[13]
port 572 nsew signal output
rlabel metal3 s 0 160080 800 160200 6 ring1_trim_a[14]
port 573 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 ring1_trim_a[15]
port 574 nsew signal output
rlabel metal3 s 0 164432 800 164552 6 ring1_trim_a[16]
port 575 nsew signal output
rlabel metal3 s 0 166472 800 166592 6 ring1_trim_a[17]
port 576 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 ring1_trim_a[18]
port 577 nsew signal output
rlabel metal3 s 0 170824 800 170944 6 ring1_trim_a[19]
port 578 nsew signal output
rlabel metal3 s 0 132064 800 132184 6 ring1_trim_a[1]
port 579 nsew signal output
rlabel metal3 s 0 173000 800 173120 6 ring1_trim_a[20]
port 580 nsew signal output
rlabel metal3 s 0 175176 800 175296 6 ring1_trim_a[21]
port 581 nsew signal output
rlabel metal3 s 0 177352 800 177472 6 ring1_trim_a[22]
port 582 nsew signal output
rlabel metal3 s 0 179392 800 179512 6 ring1_trim_a[23]
port 583 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 ring1_trim_a[24]
port 584 nsew signal output
rlabel metal3 s 0 183744 800 183864 6 ring1_trim_a[25]
port 585 nsew signal output
rlabel metal3 s 0 134240 800 134360 6 ring1_trim_a[2]
port 586 nsew signal output
rlabel metal3 s 0 136416 800 136536 6 ring1_trim_a[3]
port 587 nsew signal output
rlabel metal3 s 0 138592 800 138712 6 ring1_trim_a[4]
port 588 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 ring1_trim_a[5]
port 589 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 ring1_trim_a[6]
port 590 nsew signal output
rlabel metal3 s 0 144984 800 145104 6 ring1_trim_a[7]
port 591 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 ring1_trim_a[8]
port 592 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 ring1_trim_a[9]
port 593 nsew signal output
rlabel metal3 s 99200 189048 100000 189168 6 ring2_clk
port 594 nsew signal input
rlabel metal3 s 99200 176536 100000 176656 6 ring2_clkmux[0]
port 595 nsew signal output
rlabel metal3 s 99200 179664 100000 179784 6 ring2_clkmux[1]
port 596 nsew signal output
rlabel metal3 s 99200 182792 100000 182912 6 ring2_clkmux[2]
port 597 nsew signal output
rlabel metal3 s 99200 185920 100000 186040 6 ring2_start
port 598 nsew signal output
rlabel metal3 s 99200 1504 100000 1624 6 ring2_trim_a[0]
port 599 nsew signal output
rlabel metal3 s 99200 32648 100000 32768 6 ring2_trim_a[10]
port 600 nsew signal output
rlabel metal3 s 99200 35776 100000 35896 6 ring2_trim_a[11]
port 601 nsew signal output
rlabel metal3 s 99200 38904 100000 39024 6 ring2_trim_a[12]
port 602 nsew signal output
rlabel metal3 s 99200 42032 100000 42152 6 ring2_trim_a[13]
port 603 nsew signal output
rlabel metal3 s 99200 45160 100000 45280 6 ring2_trim_a[14]
port 604 nsew signal output
rlabel metal3 s 99200 48288 100000 48408 6 ring2_trim_a[15]
port 605 nsew signal output
rlabel metal3 s 99200 51416 100000 51536 6 ring2_trim_a[16]
port 606 nsew signal output
rlabel metal3 s 99200 54544 100000 54664 6 ring2_trim_a[17]
port 607 nsew signal output
rlabel metal3 s 99200 57672 100000 57792 6 ring2_trim_a[18]
port 608 nsew signal output
rlabel metal3 s 99200 60800 100000 60920 6 ring2_trim_a[19]
port 609 nsew signal output
rlabel metal3 s 99200 4496 100000 4616 6 ring2_trim_a[1]
port 610 nsew signal output
rlabel metal3 s 99200 63928 100000 64048 6 ring2_trim_a[20]
port 611 nsew signal output
rlabel metal3 s 99200 67056 100000 67176 6 ring2_trim_a[21]
port 612 nsew signal output
rlabel metal3 s 99200 70184 100000 70304 6 ring2_trim_a[22]
port 613 nsew signal output
rlabel metal3 s 99200 73312 100000 73432 6 ring2_trim_a[23]
port 614 nsew signal output
rlabel metal3 s 99200 76440 100000 76560 6 ring2_trim_a[24]
port 615 nsew signal output
rlabel metal3 s 99200 79568 100000 79688 6 ring2_trim_a[25]
port 616 nsew signal output
rlabel metal3 s 99200 82696 100000 82816 6 ring2_trim_a[26]
port 617 nsew signal output
rlabel metal3 s 99200 85824 100000 85944 6 ring2_trim_a[27]
port 618 nsew signal output
rlabel metal3 s 99200 7624 100000 7744 6 ring2_trim_a[2]
port 619 nsew signal output
rlabel metal3 s 99200 10752 100000 10872 6 ring2_trim_a[3]
port 620 nsew signal output
rlabel metal3 s 99200 13880 100000 14000 6 ring2_trim_a[4]
port 621 nsew signal output
rlabel metal3 s 99200 17008 100000 17128 6 ring2_trim_a[5]
port 622 nsew signal output
rlabel metal3 s 99200 20136 100000 20256 6 ring2_trim_a[6]
port 623 nsew signal output
rlabel metal3 s 99200 23264 100000 23384 6 ring2_trim_a[7]
port 624 nsew signal output
rlabel metal3 s 99200 26392 100000 26512 6 ring2_trim_a[8]
port 625 nsew signal output
rlabel metal3 s 99200 29520 100000 29640 6 ring2_trim_a[9]
port 626 nsew signal output
rlabel metal3 s 99200 88952 100000 89072 6 ring2_trim_b[0]
port 627 nsew signal output
rlabel metal3 s 99200 120232 100000 120352 6 ring2_trim_b[10]
port 628 nsew signal output
rlabel metal3 s 99200 123360 100000 123480 6 ring2_trim_b[11]
port 629 nsew signal output
rlabel metal3 s 99200 126488 100000 126608 6 ring2_trim_b[12]
port 630 nsew signal output
rlabel metal3 s 99200 129616 100000 129736 6 ring2_trim_b[13]
port 631 nsew signal output
rlabel metal3 s 99200 132744 100000 132864 6 ring2_trim_b[14]
port 632 nsew signal output
rlabel metal3 s 99200 135872 100000 135992 6 ring2_trim_b[15]
port 633 nsew signal output
rlabel metal3 s 99200 139000 100000 139120 6 ring2_trim_b[16]
port 634 nsew signal output
rlabel metal3 s 99200 142128 100000 142248 6 ring2_trim_b[17]
port 635 nsew signal output
rlabel metal3 s 99200 145256 100000 145376 6 ring2_trim_b[18]
port 636 nsew signal output
rlabel metal3 s 99200 148384 100000 148504 6 ring2_trim_b[19]
port 637 nsew signal output
rlabel metal3 s 99200 92080 100000 92200 6 ring2_trim_b[1]
port 638 nsew signal output
rlabel metal3 s 99200 151512 100000 151632 6 ring2_trim_b[20]
port 639 nsew signal output
rlabel metal3 s 99200 154640 100000 154760 6 ring2_trim_b[21]
port 640 nsew signal output
rlabel metal3 s 99200 157768 100000 157888 6 ring2_trim_b[22]
port 641 nsew signal output
rlabel metal3 s 99200 160896 100000 161016 6 ring2_trim_b[23]
port 642 nsew signal output
rlabel metal3 s 99200 164024 100000 164144 6 ring2_trim_b[24]
port 643 nsew signal output
rlabel metal3 s 99200 167152 100000 167272 6 ring2_trim_b[25]
port 644 nsew signal output
rlabel metal3 s 99200 170280 100000 170400 6 ring2_trim_b[26]
port 645 nsew signal output
rlabel metal3 s 99200 173408 100000 173528 6 ring2_trim_b[27]
port 646 nsew signal output
rlabel metal3 s 99200 95208 100000 95328 6 ring2_trim_b[2]
port 647 nsew signal output
rlabel metal3 s 99200 98336 100000 98456 6 ring2_trim_b[3]
port 648 nsew signal output
rlabel metal3 s 99200 101464 100000 101584 6 ring2_trim_b[4]
port 649 nsew signal output
rlabel metal3 s 99200 104592 100000 104712 6 ring2_trim_b[5]
port 650 nsew signal output
rlabel metal3 s 99200 107720 100000 107840 6 ring2_trim_b[6]
port 651 nsew signal output
rlabel metal3 s 99200 110848 100000 110968 6 ring2_trim_b[7]
port 652 nsew signal output
rlabel metal3 s 99200 113976 100000 114096 6 ring2_trim_b[8]
port 653 nsew signal output
rlabel metal3 s 99200 117104 100000 117224 6 ring2_trim_b[9]
port 654 nsew signal output
rlabel metal3 s 99200 192176 100000 192296 6 ring3_clk
port 655 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 ring4_clk
port 656 nsew signal input
rlabel metal3 s 0 198840 800 198960 6 ring5_clk
port 657 nsew signal input
rlabel metal3 s 99200 195304 100000 195424 6 ring6_clk
port 658 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 ring7_clk
port 659 nsew signal input
rlabel metal3 s 99200 198432 100000 198552 6 ring8_clk
port 660 nsew signal input
rlabel metal2 s 99470 199200 99526 200000 6 ring9_clk
port 661 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 662 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 663 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 663 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 663 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 664 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 665 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 666 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 667 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[10]
port 668 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[11]
port 669 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 670 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[13]
port 671 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 672 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[15]
port 673 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[16]
port 674 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[17]
port 675 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[18]
port 676 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[19]
port 677 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[1]
port 678 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[20]
port 679 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[21]
port 680 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[22]
port 681 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_adr_i[23]
port 682 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[24]
port 683 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[25]
port 684 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[26]
port 685 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[27]
port 686 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[28]
port 687 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[29]
port 688 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 689 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[30]
port 690 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[31]
port 691 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 692 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 693 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[5]
port 694 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 695 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 696 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[8]
port 697 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 698 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 699 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 700 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 701 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[11]
port 702 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 703 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[13]
port 704 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[14]
port 705 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[15]
port 706 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[16]
port 707 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 708 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[18]
port 709 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[19]
port 710 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 711 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[20]
port 712 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[21]
port 713 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[22]
port 714 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[23]
port 715 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[24]
port 716 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[25]
port 717 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[26]
port 718 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[27]
port 719 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[28]
port 720 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[29]
port 721 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[2]
port 722 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[30]
port 723 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[31]
port 724 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 725 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 726 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 727 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[6]
port 728 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 729 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[8]
port 730 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 731 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 732 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 733 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_o[11]
port 734 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[12]
port 735 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[13]
port 736 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[14]
port 737 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 738 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[16]
port 739 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[17]
port 740 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[18]
port 741 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[19]
port 742 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 743 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[20]
port 744 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[21]
port 745 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[22]
port 746 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[23]
port 747 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[24]
port 748 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[25]
port 749 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_o[26]
port 750 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[27]
port 751 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[28]
port 752 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[29]
port 753 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 754 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[30]
port 755 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_o[31]
port 756 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_o[3]
port 757 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[4]
port 758 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 759 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[6]
port 760 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 761 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 762 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[9]
port 763 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 764 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 765 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 766 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 767 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 768 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_we_i
port 769 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/digitalcore_macro/runs/digitalcore_macro/results/magic/digitalcore_macro.gds
string GDS_END 24182852
string GDS_START 764058
<< end >>

