magic
tech sky130A
magscale 1 2
timestamp 1635126048
<< obsli1 >>
rect 949 2159 98963 97393
<< obsm1 >>
rect 106 1028 99898 97708
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2962 99200 3018 100000
rect 3790 99200 3846 100000
rect 4710 99200 4766 100000
rect 5538 99200 5594 100000
rect 6458 99200 6514 100000
rect 7286 99200 7342 100000
rect 8206 99200 8262 100000
rect 9034 99200 9090 100000
rect 9862 99200 9918 100000
rect 10782 99200 10838 100000
rect 11610 99200 11666 100000
rect 12530 99200 12586 100000
rect 13358 99200 13414 100000
rect 14278 99200 14334 100000
rect 15106 99200 15162 100000
rect 16026 99200 16082 100000
rect 16854 99200 16910 100000
rect 17774 99200 17830 100000
rect 18602 99200 18658 100000
rect 19430 99200 19486 100000
rect 20350 99200 20406 100000
rect 21178 99200 21234 100000
rect 22098 99200 22154 100000
rect 22926 99200 22982 100000
rect 23846 99200 23902 100000
rect 24674 99200 24730 100000
rect 25594 99200 25650 100000
rect 26422 99200 26478 100000
rect 27342 99200 27398 100000
rect 28170 99200 28226 100000
rect 28998 99200 29054 100000
rect 29918 99200 29974 100000
rect 30746 99200 30802 100000
rect 31666 99200 31722 100000
rect 32494 99200 32550 100000
rect 33414 99200 33470 100000
rect 34242 99200 34298 100000
rect 35162 99200 35218 100000
rect 35990 99200 36046 100000
rect 36818 99200 36874 100000
rect 37738 99200 37794 100000
rect 38566 99200 38622 100000
rect 39486 99200 39542 100000
rect 40314 99200 40370 100000
rect 41234 99200 41290 100000
rect 42062 99200 42118 100000
rect 42982 99200 43038 100000
rect 43810 99200 43866 100000
rect 44730 99200 44786 100000
rect 45558 99200 45614 100000
rect 46386 99200 46442 100000
rect 47306 99200 47362 100000
rect 48134 99200 48190 100000
rect 49054 99200 49110 100000
rect 49882 99200 49938 100000
rect 50802 99200 50858 100000
rect 51630 99200 51686 100000
rect 52550 99200 52606 100000
rect 53378 99200 53434 100000
rect 54298 99200 54354 100000
rect 55126 99200 55182 100000
rect 55954 99200 56010 100000
rect 56874 99200 56930 100000
rect 57702 99200 57758 100000
rect 58622 99200 58678 100000
rect 59450 99200 59506 100000
rect 60370 99200 60426 100000
rect 61198 99200 61254 100000
rect 62118 99200 62174 100000
rect 62946 99200 63002 100000
rect 63866 99200 63922 100000
rect 64694 99200 64750 100000
rect 65522 99200 65578 100000
rect 66442 99200 66498 100000
rect 67270 99200 67326 100000
rect 68190 99200 68246 100000
rect 69018 99200 69074 100000
rect 69938 99200 69994 100000
rect 70766 99200 70822 100000
rect 71686 99200 71742 100000
rect 72514 99200 72570 100000
rect 73342 99200 73398 100000
rect 74262 99200 74318 100000
rect 75090 99200 75146 100000
rect 76010 99200 76066 100000
rect 76838 99200 76894 100000
rect 77758 99200 77814 100000
rect 78586 99200 78642 100000
rect 79506 99200 79562 100000
rect 80334 99200 80390 100000
rect 81254 99200 81310 100000
rect 82082 99200 82138 100000
rect 82910 99200 82966 100000
rect 83830 99200 83886 100000
rect 84658 99200 84714 100000
rect 85578 99200 85634 100000
rect 86406 99200 86462 100000
rect 87326 99200 87382 100000
rect 88154 99200 88210 100000
rect 89074 99200 89130 100000
rect 89902 99200 89958 100000
rect 90822 99200 90878 100000
rect 91650 99200 91706 100000
rect 92478 99200 92534 100000
rect 93398 99200 93454 100000
rect 94226 99200 94282 100000
rect 95146 99200 95202 100000
rect 95974 99200 96030 100000
rect 96894 99200 96950 100000
rect 97722 99200 97778 100000
rect 98642 99200 98698 100000
rect 99470 99200 99526 100000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62946 0 63002 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72882 0 72938 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82634 0 82690 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 112 99144 330 99385
rect 498 99144 1158 99385
rect 1326 99144 1986 99385
rect 2154 99144 2906 99385
rect 3074 99144 3734 99385
rect 3902 99144 4654 99385
rect 4822 99144 5482 99385
rect 5650 99144 6402 99385
rect 6570 99144 7230 99385
rect 7398 99144 8150 99385
rect 8318 99144 8978 99385
rect 9146 99144 9806 99385
rect 9974 99144 10726 99385
rect 10894 99144 11554 99385
rect 11722 99144 12474 99385
rect 12642 99144 13302 99385
rect 13470 99144 14222 99385
rect 14390 99144 15050 99385
rect 15218 99144 15970 99385
rect 16138 99144 16798 99385
rect 16966 99144 17718 99385
rect 17886 99144 18546 99385
rect 18714 99144 19374 99385
rect 19542 99144 20294 99385
rect 20462 99144 21122 99385
rect 21290 99144 22042 99385
rect 22210 99144 22870 99385
rect 23038 99144 23790 99385
rect 23958 99144 24618 99385
rect 24786 99144 25538 99385
rect 25706 99144 26366 99385
rect 26534 99144 27286 99385
rect 27454 99144 28114 99385
rect 28282 99144 28942 99385
rect 29110 99144 29862 99385
rect 30030 99144 30690 99385
rect 30858 99144 31610 99385
rect 31778 99144 32438 99385
rect 32606 99144 33358 99385
rect 33526 99144 34186 99385
rect 34354 99144 35106 99385
rect 35274 99144 35934 99385
rect 36102 99144 36762 99385
rect 36930 99144 37682 99385
rect 37850 99144 38510 99385
rect 38678 99144 39430 99385
rect 39598 99144 40258 99385
rect 40426 99144 41178 99385
rect 41346 99144 42006 99385
rect 42174 99144 42926 99385
rect 43094 99144 43754 99385
rect 43922 99144 44674 99385
rect 44842 99144 45502 99385
rect 45670 99144 46330 99385
rect 46498 99144 47250 99385
rect 47418 99144 48078 99385
rect 48246 99144 48998 99385
rect 49166 99144 49826 99385
rect 49994 99144 50746 99385
rect 50914 99144 51574 99385
rect 51742 99144 52494 99385
rect 52662 99144 53322 99385
rect 53490 99144 54242 99385
rect 54410 99144 55070 99385
rect 55238 99144 55898 99385
rect 56066 99144 56818 99385
rect 56986 99144 57646 99385
rect 57814 99144 58566 99385
rect 58734 99144 59394 99385
rect 59562 99144 60314 99385
rect 60482 99144 61142 99385
rect 61310 99144 62062 99385
rect 62230 99144 62890 99385
rect 63058 99144 63810 99385
rect 63978 99144 64638 99385
rect 64806 99144 65466 99385
rect 65634 99144 66386 99385
rect 66554 99144 67214 99385
rect 67382 99144 68134 99385
rect 68302 99144 68962 99385
rect 69130 99144 69882 99385
rect 70050 99144 70710 99385
rect 70878 99144 71630 99385
rect 71798 99144 72458 99385
rect 72626 99144 73286 99385
rect 73454 99144 74206 99385
rect 74374 99144 75034 99385
rect 75202 99144 75954 99385
rect 76122 99144 76782 99385
rect 76950 99144 77702 99385
rect 77870 99144 78530 99385
rect 78698 99144 79450 99385
rect 79618 99144 80278 99385
rect 80446 99144 81198 99385
rect 81366 99144 82026 99385
rect 82194 99144 82854 99385
rect 83022 99144 83774 99385
rect 83942 99144 84602 99385
rect 84770 99144 85522 99385
rect 85690 99144 86350 99385
rect 86518 99144 87270 99385
rect 87438 99144 88098 99385
rect 88266 99144 89018 99385
rect 89186 99144 89846 99385
rect 90014 99144 90766 99385
rect 90934 99144 91594 99385
rect 91762 99144 92422 99385
rect 92590 99144 93342 99385
rect 93510 99144 94170 99385
rect 94338 99144 95090 99385
rect 95258 99144 95918 99385
rect 96086 99144 96838 99385
rect 97006 99144 97666 99385
rect 97834 99144 98586 99385
rect 98754 99144 99414 99385
rect 99582 99144 99892 99385
rect 112 856 99892 99144
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 606 856
rect 774 800 790 856
rect 958 800 1066 856
rect 1234 800 1250 856
rect 1418 800 1434 856
rect 1602 800 1618 856
rect 1786 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2262 856
rect 2430 800 2446 856
rect 2614 800 2630 856
rect 2798 800 2814 856
rect 2982 800 3090 856
rect 3258 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3826 856
rect 3994 800 4102 856
rect 4270 800 4286 856
rect 4454 800 4470 856
rect 4638 800 4654 856
rect 4822 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5666 856
rect 5834 800 5850 856
rect 6018 800 6126 856
rect 6294 800 6310 856
rect 6478 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7690 856
rect 7858 800 7874 856
rect 8042 800 8150 856
rect 8318 800 8334 856
rect 8502 800 8518 856
rect 8686 800 8702 856
rect 8870 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9346 856
rect 9514 800 9530 856
rect 9698 800 9714 856
rect 9882 800 9990 856
rect 10158 800 10174 856
rect 10342 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10726 856
rect 10894 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11554 856
rect 11722 800 11738 856
rect 11906 800 12014 856
rect 12182 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12566 856
rect 12734 800 12750 856
rect 12918 800 13026 856
rect 13194 800 13210 856
rect 13378 800 13394 856
rect 13562 800 13578 856
rect 13746 800 13762 856
rect 13930 800 14038 856
rect 14206 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14590 856
rect 14758 800 14774 856
rect 14942 800 15050 856
rect 15218 800 15234 856
rect 15402 800 15418 856
rect 15586 800 15602 856
rect 15770 800 15786 856
rect 15954 800 16062 856
rect 16230 800 16246 856
rect 16414 800 16430 856
rect 16598 800 16614 856
rect 16782 800 16890 856
rect 17058 800 17074 856
rect 17242 800 17258 856
rect 17426 800 17442 856
rect 17610 800 17626 856
rect 17794 800 17902 856
rect 18070 800 18086 856
rect 18254 800 18270 856
rect 18438 800 18454 856
rect 18622 800 18638 856
rect 18806 800 18914 856
rect 19082 800 19098 856
rect 19266 800 19282 856
rect 19450 800 19466 856
rect 19634 800 19650 856
rect 19818 800 19926 856
rect 20094 800 20110 856
rect 20278 800 20294 856
rect 20462 800 20478 856
rect 20646 800 20662 856
rect 20830 800 20938 856
rect 21106 800 21122 856
rect 21290 800 21306 856
rect 21474 800 21490 856
rect 21658 800 21674 856
rect 21842 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22318 856
rect 22486 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22962 856
rect 23130 800 23146 856
rect 23314 800 23330 856
rect 23498 800 23514 856
rect 23682 800 23698 856
rect 23866 800 23974 856
rect 24142 800 24158 856
rect 24326 800 24342 856
rect 24510 800 24526 856
rect 24694 800 24710 856
rect 24878 800 24986 856
rect 25154 800 25170 856
rect 25338 800 25354 856
rect 25522 800 25538 856
rect 25706 800 25814 856
rect 25982 800 25998 856
rect 26166 800 26182 856
rect 26350 800 26366 856
rect 26534 800 26550 856
rect 26718 800 26826 856
rect 26994 800 27010 856
rect 27178 800 27194 856
rect 27362 800 27378 856
rect 27546 800 27562 856
rect 27730 800 27838 856
rect 28006 800 28022 856
rect 28190 800 28206 856
rect 28374 800 28390 856
rect 28558 800 28574 856
rect 28742 800 28850 856
rect 29018 800 29034 856
rect 29202 800 29218 856
rect 29386 800 29402 856
rect 29570 800 29586 856
rect 29754 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30230 856
rect 30398 800 30414 856
rect 30582 800 30598 856
rect 30766 800 30874 856
rect 31042 800 31058 856
rect 31226 800 31242 856
rect 31410 800 31426 856
rect 31594 800 31610 856
rect 31778 800 31886 856
rect 32054 800 32070 856
rect 32238 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33266 856
rect 33434 800 33450 856
rect 33618 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34094 856
rect 34262 800 34278 856
rect 34446 800 34462 856
rect 34630 800 34738 856
rect 34906 800 34922 856
rect 35090 800 35106 856
rect 35274 800 35290 856
rect 35458 800 35474 856
rect 35642 800 35750 856
rect 35918 800 35934 856
rect 36102 800 36118 856
rect 36286 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36762 856
rect 36930 800 36946 856
rect 37114 800 37130 856
rect 37298 800 37314 856
rect 37482 800 37498 856
rect 37666 800 37774 856
rect 37942 800 37958 856
rect 38126 800 38142 856
rect 38310 800 38326 856
rect 38494 800 38510 856
rect 38678 800 38786 856
rect 38954 800 38970 856
rect 39138 800 39154 856
rect 39322 800 39338 856
rect 39506 800 39522 856
rect 39690 800 39798 856
rect 39966 800 39982 856
rect 40150 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40534 856
rect 40702 800 40810 856
rect 40978 800 40994 856
rect 41162 800 41178 856
rect 41346 800 41362 856
rect 41530 800 41546 856
rect 41714 800 41822 856
rect 41990 800 42006 856
rect 42174 800 42190 856
rect 42358 800 42374 856
rect 42542 800 42650 856
rect 42818 800 42834 856
rect 43002 800 43018 856
rect 43186 800 43202 856
rect 43370 800 43386 856
rect 43554 800 43662 856
rect 43830 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44398 856
rect 44566 800 44674 856
rect 44842 800 44858 856
rect 45026 800 45042 856
rect 45210 800 45226 856
rect 45394 800 45410 856
rect 45578 800 45686 856
rect 45854 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46238 856
rect 46406 800 46422 856
rect 46590 800 46698 856
rect 46866 800 46882 856
rect 47050 800 47066 856
rect 47234 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48262 856
rect 48430 800 48446 856
rect 48614 800 48722 856
rect 48890 800 48906 856
rect 49074 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49458 856
rect 49626 800 49734 856
rect 49902 800 49918 856
rect 50086 800 50102 856
rect 50270 800 50286 856
rect 50454 800 50562 856
rect 50730 800 50746 856
rect 50914 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51298 856
rect 51466 800 51574 856
rect 51742 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52126 856
rect 52294 800 52310 856
rect 52478 800 52586 856
rect 52754 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53138 856
rect 53306 800 53322 856
rect 53490 800 53598 856
rect 53766 800 53782 856
rect 53950 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54334 856
rect 54502 800 54610 856
rect 54778 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55162 856
rect 55330 800 55346 856
rect 55514 800 55622 856
rect 55790 800 55806 856
rect 55974 800 55990 856
rect 56158 800 56174 856
rect 56342 800 56358 856
rect 56526 800 56634 856
rect 56802 800 56818 856
rect 56986 800 57002 856
rect 57170 800 57186 856
rect 57354 800 57370 856
rect 57538 800 57646 856
rect 57814 800 57830 856
rect 57998 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58842 856
rect 59010 800 59026 856
rect 59194 800 59210 856
rect 59378 800 59486 856
rect 59654 800 59670 856
rect 59838 800 59854 856
rect 60022 800 60038 856
rect 60206 800 60222 856
rect 60390 800 60498 856
rect 60666 800 60682 856
rect 60850 800 60866 856
rect 61034 800 61050 856
rect 61218 800 61234 856
rect 61402 800 61510 856
rect 61678 800 61694 856
rect 61862 800 61878 856
rect 62046 800 62062 856
rect 62230 800 62246 856
rect 62414 800 62522 856
rect 62690 800 62706 856
rect 62874 800 62890 856
rect 63058 800 63074 856
rect 63242 800 63258 856
rect 63426 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63902 856
rect 64070 800 64086 856
rect 64254 800 64270 856
rect 64438 800 64546 856
rect 64714 800 64730 856
rect 64898 800 64914 856
rect 65082 800 65098 856
rect 65266 800 65282 856
rect 65450 800 65558 856
rect 65726 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66110 856
rect 66278 800 66294 856
rect 66462 800 66570 856
rect 66738 800 66754 856
rect 66922 800 66938 856
rect 67106 800 67122 856
rect 67290 800 67398 856
rect 67566 800 67582 856
rect 67750 800 67766 856
rect 67934 800 67950 856
rect 68118 800 68134 856
rect 68302 800 68410 856
rect 68578 800 68594 856
rect 68762 800 68778 856
rect 68946 800 68962 856
rect 69130 800 69146 856
rect 69314 800 69422 856
rect 69590 800 69606 856
rect 69774 800 69790 856
rect 69958 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70434 856
rect 70602 800 70618 856
rect 70786 800 70802 856
rect 70970 800 70986 856
rect 71154 800 71170 856
rect 71338 800 71446 856
rect 71614 800 71630 856
rect 71798 800 71814 856
rect 71982 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72458 856
rect 72626 800 72642 856
rect 72810 800 72826 856
rect 72994 800 73010 856
rect 73178 800 73194 856
rect 73362 800 73470 856
rect 73638 800 73654 856
rect 73822 800 73838 856
rect 74006 800 74022 856
rect 74190 800 74206 856
rect 74374 800 74482 856
rect 74650 800 74666 856
rect 74834 800 74850 856
rect 75018 800 75034 856
rect 75202 800 75310 856
rect 75478 800 75494 856
rect 75662 800 75678 856
rect 75846 800 75862 856
rect 76030 800 76046 856
rect 76214 800 76322 856
rect 76490 800 76506 856
rect 76674 800 76690 856
rect 76858 800 76874 856
rect 77042 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77518 856
rect 77686 800 77702 856
rect 77870 800 77886 856
rect 78054 800 78070 856
rect 78238 800 78346 856
rect 78514 800 78530 856
rect 78698 800 78714 856
rect 78882 800 78898 856
rect 79066 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79726 856
rect 79894 800 79910 856
rect 80078 800 80094 856
rect 80262 800 80370 856
rect 80538 800 80554 856
rect 80722 800 80738 856
rect 80906 800 80922 856
rect 81090 800 81106 856
rect 81274 800 81382 856
rect 81550 800 81566 856
rect 81734 800 81750 856
rect 81918 800 81934 856
rect 82102 800 82118 856
rect 82286 800 82394 856
rect 82562 800 82578 856
rect 82746 800 82762 856
rect 82930 800 82946 856
rect 83114 800 83130 856
rect 83298 800 83406 856
rect 83574 800 83590 856
rect 83758 800 83774 856
rect 83942 800 83958 856
rect 84126 800 84234 856
rect 84402 800 84418 856
rect 84586 800 84602 856
rect 84770 800 84786 856
rect 84954 800 84970 856
rect 85138 800 85246 856
rect 85414 800 85430 856
rect 85598 800 85614 856
rect 85782 800 85798 856
rect 85966 800 85982 856
rect 86150 800 86258 856
rect 86426 800 86442 856
rect 86610 800 86626 856
rect 86794 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87270 856
rect 87438 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88006 856
rect 88174 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88650 856
rect 88818 800 88834 856
rect 89002 800 89018 856
rect 89186 800 89294 856
rect 89462 800 89478 856
rect 89646 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90030 856
rect 90198 800 90306 856
rect 90474 800 90490 856
rect 90658 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91042 856
rect 91210 800 91318 856
rect 91486 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91870 856
rect 92038 800 92146 856
rect 92314 800 92330 856
rect 92498 800 92514 856
rect 92682 800 92698 856
rect 92866 800 92882 856
rect 93050 800 93158 856
rect 93326 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93710 856
rect 93878 800 93894 856
rect 94062 800 94170 856
rect 94338 800 94354 856
rect 94522 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95734 856
rect 95902 800 95918 856
rect 96086 800 96194 856
rect 96362 800 96378 856
rect 96546 800 96562 856
rect 96730 800 96746 856
rect 96914 800 96930 856
rect 97098 800 97206 856
rect 97374 800 97390 856
rect 97558 800 97574 856
rect 97742 800 97758 856
rect 97926 800 97942 856
rect 98110 800 98218 856
rect 98386 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 98954 856
rect 99122 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99598 856
rect 99766 800 99782 856
<< metal3 >>
rect 0 99288 800 99408
rect 0 98200 800 98320
rect 0 97112 800 97232
rect 0 96024 800 96144
rect 0 94936 800 95056
rect 0 93848 800 93968
rect 0 92760 800 92880
rect 0 91672 800 91792
rect 0 90584 800 90704
rect 0 89496 800 89616
rect 0 88408 800 88528
rect 0 87320 800 87440
rect 0 86232 800 86352
rect 0 85008 800 85128
rect 0 83920 800 84040
rect 0 82832 800 82952
rect 0 81744 800 81864
rect 0 80656 800 80776
rect 0 79568 800 79688
rect 0 78480 800 78600
rect 0 77392 800 77512
rect 0 76304 800 76424
rect 0 75216 800 75336
rect 0 74128 800 74248
rect 0 73040 800 73160
rect 0 71952 800 72072
rect 0 70728 800 70848
rect 0 69640 800 69760
rect 0 68552 800 68672
rect 0 67464 800 67584
rect 0 66376 800 66496
rect 0 65288 800 65408
rect 0 64200 800 64320
rect 0 63112 800 63232
rect 0 62024 800 62144
rect 0 60936 800 61056
rect 0 59848 800 59968
rect 0 58760 800 58880
rect 0 57672 800 57792
rect 0 56448 800 56568
rect 0 55360 800 55480
rect 0 54272 800 54392
rect 0 53184 800 53304
rect 0 52096 800 52216
rect 0 51008 800 51128
rect 0 49920 800 50040
rect 0 48832 800 48952
rect 0 47744 800 47864
rect 0 46656 800 46776
rect 0 45568 800 45688
rect 0 44480 800 44600
rect 0 43392 800 43512
rect 0 42168 800 42288
rect 0 41080 800 41200
rect 0 39992 800 40112
rect 0 38904 800 39024
rect 0 37816 800 37936
rect 0 36728 800 36848
rect 0 35640 800 35760
rect 0 34552 800 34672
rect 0 33464 800 33584
rect 0 32376 800 32496
rect 0 31288 800 31408
rect 0 30200 800 30320
rect 0 29112 800 29232
rect 0 27888 800 28008
rect 0 26800 800 26920
rect 0 25712 800 25832
rect 0 24624 800 24744
rect 0 23536 800 23656
rect 0 22448 800 22568
rect 0 21360 800 21480
rect 0 20272 800 20392
rect 0 19184 800 19304
rect 0 18096 800 18216
rect 0 17008 800 17128
rect 0 15920 800 16040
rect 0 14832 800 14952
rect 0 13608 800 13728
rect 0 12520 800 12640
rect 0 11432 800 11552
rect 0 10344 800 10464
rect 0 9256 800 9376
rect 0 8168 800 8288
rect 0 7080 800 7200
rect 0 5992 800 6112
rect 0 4904 800 5024
rect 0 3816 800 3936
rect 0 2728 800 2848
rect 0 1640 800 1760
rect 0 552 800 672
<< obsm3 >>
rect 880 99208 97875 99381
rect 381 98400 97875 99208
rect 880 98120 97875 98400
rect 381 97312 97875 98120
rect 880 97032 97875 97312
rect 381 96224 97875 97032
rect 880 95944 97875 96224
rect 381 95136 97875 95944
rect 880 94856 97875 95136
rect 381 94048 97875 94856
rect 880 93768 97875 94048
rect 381 92960 97875 93768
rect 880 92680 97875 92960
rect 381 91872 97875 92680
rect 880 91592 97875 91872
rect 381 90784 97875 91592
rect 880 90504 97875 90784
rect 381 89696 97875 90504
rect 880 89416 97875 89696
rect 381 88608 97875 89416
rect 880 88328 97875 88608
rect 381 87520 97875 88328
rect 880 87240 97875 87520
rect 381 86432 97875 87240
rect 880 86152 97875 86432
rect 381 85208 97875 86152
rect 880 84928 97875 85208
rect 381 84120 97875 84928
rect 880 83840 97875 84120
rect 381 83032 97875 83840
rect 880 82752 97875 83032
rect 381 81944 97875 82752
rect 880 81664 97875 81944
rect 381 80856 97875 81664
rect 880 80576 97875 80856
rect 381 79768 97875 80576
rect 880 79488 97875 79768
rect 381 78680 97875 79488
rect 880 78400 97875 78680
rect 381 77592 97875 78400
rect 880 77312 97875 77592
rect 381 76504 97875 77312
rect 880 76224 97875 76504
rect 381 75416 97875 76224
rect 880 75136 97875 75416
rect 381 74328 97875 75136
rect 880 74048 97875 74328
rect 381 73240 97875 74048
rect 880 72960 97875 73240
rect 381 72152 97875 72960
rect 880 71872 97875 72152
rect 381 70928 97875 71872
rect 880 70648 97875 70928
rect 381 69840 97875 70648
rect 880 69560 97875 69840
rect 381 68752 97875 69560
rect 880 68472 97875 68752
rect 381 67664 97875 68472
rect 880 67384 97875 67664
rect 381 66576 97875 67384
rect 880 66296 97875 66576
rect 381 65488 97875 66296
rect 880 65208 97875 65488
rect 381 64400 97875 65208
rect 880 64120 97875 64400
rect 381 63312 97875 64120
rect 880 63032 97875 63312
rect 381 62224 97875 63032
rect 880 61944 97875 62224
rect 381 61136 97875 61944
rect 880 60856 97875 61136
rect 381 60048 97875 60856
rect 880 59768 97875 60048
rect 381 58960 97875 59768
rect 880 58680 97875 58960
rect 381 57872 97875 58680
rect 880 57592 97875 57872
rect 381 56648 97875 57592
rect 880 56368 97875 56648
rect 381 55560 97875 56368
rect 880 55280 97875 55560
rect 381 54472 97875 55280
rect 880 54192 97875 54472
rect 381 53384 97875 54192
rect 880 53104 97875 53384
rect 381 52296 97875 53104
rect 880 52016 97875 52296
rect 381 51208 97875 52016
rect 880 50928 97875 51208
rect 381 50120 97875 50928
rect 880 49840 97875 50120
rect 381 49032 97875 49840
rect 880 48752 97875 49032
rect 381 47944 97875 48752
rect 880 47664 97875 47944
rect 381 46856 97875 47664
rect 880 46576 97875 46856
rect 381 45768 97875 46576
rect 880 45488 97875 45768
rect 381 44680 97875 45488
rect 880 44400 97875 44680
rect 381 43592 97875 44400
rect 880 43312 97875 43592
rect 381 42368 97875 43312
rect 880 42088 97875 42368
rect 381 41280 97875 42088
rect 880 41000 97875 41280
rect 381 40192 97875 41000
rect 880 39912 97875 40192
rect 381 39104 97875 39912
rect 880 38824 97875 39104
rect 381 38016 97875 38824
rect 880 37736 97875 38016
rect 381 36928 97875 37736
rect 880 36648 97875 36928
rect 381 35840 97875 36648
rect 880 35560 97875 35840
rect 381 34752 97875 35560
rect 880 34472 97875 34752
rect 381 33664 97875 34472
rect 880 33384 97875 33664
rect 381 32576 97875 33384
rect 880 32296 97875 32576
rect 381 31488 97875 32296
rect 880 31208 97875 31488
rect 381 30400 97875 31208
rect 880 30120 97875 30400
rect 381 29312 97875 30120
rect 880 29032 97875 29312
rect 381 28088 97875 29032
rect 880 27808 97875 28088
rect 381 27000 97875 27808
rect 880 26720 97875 27000
rect 381 25912 97875 26720
rect 880 25632 97875 25912
rect 381 24824 97875 25632
rect 880 24544 97875 24824
rect 381 23736 97875 24544
rect 880 23456 97875 23736
rect 381 22648 97875 23456
rect 880 22368 97875 22648
rect 381 21560 97875 22368
rect 880 21280 97875 21560
rect 381 20472 97875 21280
rect 880 20192 97875 20472
rect 381 19384 97875 20192
rect 880 19104 97875 19384
rect 381 18296 97875 19104
rect 880 18016 97875 18296
rect 381 17208 97875 18016
rect 880 16928 97875 17208
rect 381 16120 97875 16928
rect 880 15840 97875 16120
rect 381 15032 97875 15840
rect 880 14752 97875 15032
rect 381 13808 97875 14752
rect 880 13528 97875 13808
rect 381 12720 97875 13528
rect 880 12440 97875 12720
rect 381 11632 97875 12440
rect 880 11352 97875 11632
rect 381 10544 97875 11352
rect 880 10264 97875 10544
rect 381 9456 97875 10264
rect 880 9176 97875 9456
rect 381 8368 97875 9176
rect 880 8088 97875 8368
rect 381 7280 97875 8088
rect 880 7000 97875 7280
rect 381 6192 97875 7000
rect 880 5912 97875 6192
rect 381 5104 97875 5912
rect 880 4824 97875 5104
rect 381 4016 97875 4824
rect 880 3736 97875 4016
rect 381 2928 97875 3736
rect 880 2648 97875 2928
rect 381 1840 97875 2648
rect 880 1560 97875 1840
rect 381 752 97875 1560
rect 880 582 97875 752
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 979 2048 4128 95573
rect 4608 2048 19488 95573
rect 19968 2048 34848 95573
rect 35328 2048 49437 95573
rect 979 987 49437 2048
<< labels >>
rlabel metal2 s 386 99200 442 100000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26422 99200 26478 100000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 28998 99200 29054 100000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31666 99200 31722 100000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34242 99200 34298 100000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 36818 99200 36874 100000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39486 99200 39542 100000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42062 99200 42118 100000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 44730 99200 44786 100000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47306 99200 47362 100000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 49882 99200 49938 100000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 99200 3018 100000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 52550 99200 52606 100000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55126 99200 55182 100000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57702 99200 57758 100000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60370 99200 60426 100000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 62946 99200 63002 100000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 65522 99200 65578 100000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70766 99200 70822 100000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73342 99200 73398 100000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76010 99200 76066 100000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5538 99200 5594 100000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81254 99200 81310 100000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 83830 99200 83886 100000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 86406 99200 86462 100000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89074 99200 89130 100000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 91650 99200 91706 100000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 94226 99200 94282 100000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 96894 99200 96950 100000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 99200 8262 100000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10782 99200 10838 100000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13358 99200 13414 100000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16026 99200 16082 100000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18602 99200 18658 100000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21178 99200 21234 100000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23846 99200 23902 100000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27342 99200 27398 100000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 29918 99200 29974 100000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32494 99200 32550 100000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35162 99200 35218 100000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 37738 99200 37794 100000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40314 99200 40370 100000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 42982 99200 43038 100000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45558 99200 45614 100000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48134 99200 48190 100000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 50802 99200 50858 100000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3790 99200 3846 100000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53378 99200 53434 100000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 55954 99200 56010 100000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 58622 99200 58678 100000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61198 99200 61254 100000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 63866 99200 63922 100000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66442 99200 66498 100000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69018 99200 69074 100000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 71686 99200 71742 100000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74262 99200 74318 100000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 76838 99200 76894 100000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 99200 6514 100000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 79506 99200 79562 100000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82082 99200 82138 100000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 84658 99200 84714 100000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 87326 99200 87382 100000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 89902 99200 89958 100000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 92478 99200 92534 100000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95146 99200 95202 100000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 97722 99200 97778 100000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9034 99200 9090 100000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11610 99200 11666 100000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14278 99200 14334 100000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 16854 99200 16910 100000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19430 99200 19486 100000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22098 99200 22154 100000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24674 99200 24730 100000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2042 99200 2098 100000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28170 99200 28226 100000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 30746 99200 30802 100000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33414 99200 33470 100000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 35990 99200 36046 100000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38566 99200 38622 100000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41234 99200 41290 100000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 43810 99200 43866 100000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46386 99200 46442 100000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49054 99200 49110 100000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 51630 99200 51686 100000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54298 99200 54354 100000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 56874 99200 56930 100000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 59450 99200 59506 100000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62118 99200 62174 100000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 64694 99200 64750 100000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67270 99200 67326 100000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 69938 99200 69994 100000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 72514 99200 72570 100000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75090 99200 75146 100000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 77758 99200 77814 100000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7286 99200 7342 100000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 80334 99200 80390 100000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 82910 99200 82966 100000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 85578 99200 85634 100000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88154 99200 88210 100000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 90822 99200 90878 100000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 93398 99200 93454 100000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 98642 99200 98698 100000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9862 99200 9918 100000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12530 99200 12586 100000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15106 99200 15162 100000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17774 99200 17830 100000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20350 99200 20406 100000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22926 99200 22982 100000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25594 99200 25650 100000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 99470 99200 99526 100000 6 ring0_clk
port 502 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 ring0_clkmux[0]
port 503 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 ring0_clkmux[1]
port 504 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 ring0_clkmux[2]
port 505 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 ring0_start
port 506 nsew signal output
rlabel metal3 s 0 552 800 672 6 ring0_trim_a[0]
port 507 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 ring0_trim_a[10]
port 508 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 ring0_trim_a[11]
port 509 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 ring0_trim_a[12]
port 510 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 ring0_trim_a[13]
port 511 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 ring0_trim_a[14]
port 512 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 ring0_trim_a[15]
port 513 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 ring0_trim_a[16]
port 514 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 ring0_trim_a[17]
port 515 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 ring0_trim_a[18]
port 516 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 ring0_trim_a[19]
port 517 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 ring0_trim_a[1]
port 518 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 ring0_trim_a[20]
port 519 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 ring0_trim_a[21]
port 520 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 ring0_trim_a[22]
port 521 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 ring0_trim_a[23]
port 522 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 ring0_trim_a[24]
port 523 nsew signal output
rlabel metal3 s 0 55360 800 55480 6 ring0_trim_a[25]
port 524 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 ring0_trim_a[26]
port 525 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 ring0_trim_a[27]
port 526 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 ring0_trim_a[2]
port 527 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 ring0_trim_a[3]
port 528 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 ring0_trim_a[4]
port 529 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 ring0_trim_a[5]
port 530 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 ring0_trim_a[6]
port 531 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 ring0_trim_a[7]
port 532 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 ring0_trim_a[8]
port 533 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 ring0_trim_a[9]
port 534 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 ring0_trim_b[0]
port 535 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 ring0_trim_b[10]
port 536 nsew signal output
rlabel metal3 s 0 71952 800 72072 6 ring0_trim_b[11]
port 537 nsew signal output
rlabel metal3 s 0 73040 800 73160 6 ring0_trim_b[12]
port 538 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 ring0_trim_b[13]
port 539 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 ring0_trim_b[14]
port 540 nsew signal output
rlabel metal3 s 0 76304 800 76424 6 ring0_trim_b[15]
port 541 nsew signal output
rlabel metal3 s 0 77392 800 77512 6 ring0_trim_b[16]
port 542 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 ring0_trim_b[17]
port 543 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 ring0_trim_b[18]
port 544 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 ring0_trim_b[19]
port 545 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 ring0_trim_b[1]
port 546 nsew signal output
rlabel metal3 s 0 81744 800 81864 6 ring0_trim_b[20]
port 547 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 ring0_trim_b[21]
port 548 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 ring0_trim_b[22]
port 549 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 ring0_trim_b[23]
port 550 nsew signal output
rlabel metal3 s 0 86232 800 86352 6 ring0_trim_b[24]
port 551 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 ring0_trim_b[25]
port 552 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 ring0_trim_b[26]
port 553 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 ring0_trim_b[27]
port 554 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 ring0_trim_b[2]
port 555 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 ring0_trim_b[3]
port 556 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 ring0_trim_b[4]
port 557 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 ring0_trim_b[5]
port 558 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 ring0_trim_b[6]
port 559 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 ring0_trim_b[7]
port 560 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 ring0_trim_b[8]
port 561 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 ring0_trim_b[9]
port 562 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 ring1_clk
port 563 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 ring1_clkmux[0]
port 564 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 ring1_clkmux[1]
port 565 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 ring1_clkmux[2]
port 566 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 ring1_start
port 567 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 ring1_trim_a[0]
port 568 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 ring1_trim_a[10]
port 569 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 ring1_trim_a[11]
port 570 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 ring1_trim_a[12]
port 571 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 ring1_trim_a[13]
port 572 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 ring1_trim_a[14]
port 573 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 ring1_trim_a[15]
port 574 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 ring1_trim_a[16]
port 575 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 ring1_trim_a[17]
port 576 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 ring1_trim_a[18]
port 577 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 ring1_trim_a[19]
port 578 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 ring1_trim_a[1]
port 579 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 ring1_trim_a[20]
port 580 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 ring1_trim_a[21]
port 581 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 ring1_trim_a[22]
port 582 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 ring1_trim_a[23]
port 583 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 ring1_trim_a[24]
port 584 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 ring1_trim_a[25]
port 585 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 ring1_trim_a[2]
port 586 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 ring1_trim_a[3]
port 587 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 ring1_trim_a[4]
port 588 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 ring1_trim_a[5]
port 589 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 ring1_trim_a[6]
port 590 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 ring1_trim_a[7]
port 591 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 ring1_trim_a[8]
port 592 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 ring1_trim_a[9]
port 593 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 595 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 595 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 595 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 596 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 597 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 598 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 599 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 600 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[11]
port 601 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 602 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 603 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 604 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 605 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[16]
port 606 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 607 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 608 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[19]
port 609 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 610 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 611 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[21]
port 612 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 613 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 614 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[24]
port 615 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 616 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 617 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[27]
port 618 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[28]
port 619 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[29]
port 620 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 621 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 622 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[31]
port 623 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 624 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 625 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 626 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 627 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 628 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[8]
port 629 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 630 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 631 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 632 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 633 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 634 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 635 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 636 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[14]
port 637 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 638 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 639 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 640 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 641 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[19]
port 642 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 643 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 644 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 645 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[22]
port 646 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 647 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 648 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[25]
port 649 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[26]
port 650 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[27]
port 651 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 652 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 653 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 654 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[30]
port 655 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[31]
port 656 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 657 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 658 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 659 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[6]
port 660 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 661 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 662 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 663 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 664 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 665 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 666 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[12]
port 667 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 668 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 669 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 670 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 671 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[17]
port 672 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 673 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 674 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 675 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[20]
port 676 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 677 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[22]
port 678 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 679 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 680 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[25]
port 681 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 682 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 683 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[28]
port 684 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[29]
port 685 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 686 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[30]
port 687 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 688 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 689 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[4]
port 690 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 691 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 692 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 693 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 694 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[9]
port 695 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 696 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 697 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 698 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 699 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 700 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 701 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 100000
string LEFview TRUE
string GDS_FILE /project/openlane/digitalcore_macro/runs/digitalcore_macro/results/magic/digitalcore_macro.gds
string GDS_END 12567730
string GDS_START 706646
<< end >>

