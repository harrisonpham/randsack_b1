magic
tech sky130A
magscale 1 2
timestamp 1635318596
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 1028 99898 97640
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2134 99200 2190 100000
rect 2962 99200 3018 100000
rect 3882 99200 3938 100000
rect 4710 99200 4766 100000
rect 5630 99200 5686 100000
rect 6458 99200 6514 100000
rect 7378 99200 7434 100000
rect 8206 99200 8262 100000
rect 9126 99200 9182 100000
rect 9954 99200 10010 100000
rect 10874 99200 10930 100000
rect 11702 99200 11758 100000
rect 12622 99200 12678 100000
rect 13542 99200 13598 100000
rect 14370 99200 14426 100000
rect 15290 99200 15346 100000
rect 16118 99200 16174 100000
rect 17038 99200 17094 100000
rect 17866 99200 17922 100000
rect 18786 99200 18842 100000
rect 19614 99200 19670 100000
rect 20534 99200 20590 100000
rect 21362 99200 21418 100000
rect 22282 99200 22338 100000
rect 23110 99200 23166 100000
rect 24030 99200 24086 100000
rect 24858 99200 24914 100000
rect 25778 99200 25834 100000
rect 26698 99200 26754 100000
rect 27526 99200 27582 100000
rect 28446 99200 28502 100000
rect 29274 99200 29330 100000
rect 30194 99200 30250 100000
rect 31022 99200 31078 100000
rect 31942 99200 31998 100000
rect 32770 99200 32826 100000
rect 33690 99200 33746 100000
rect 34518 99200 34574 100000
rect 35438 99200 35494 100000
rect 36266 99200 36322 100000
rect 37186 99200 37242 100000
rect 38106 99200 38162 100000
rect 38934 99200 38990 100000
rect 39854 99200 39910 100000
rect 40682 99200 40738 100000
rect 41602 99200 41658 100000
rect 42430 99200 42486 100000
rect 43350 99200 43406 100000
rect 44178 99200 44234 100000
rect 45098 99200 45154 100000
rect 45926 99200 45982 100000
rect 46846 99200 46902 100000
rect 47674 99200 47730 100000
rect 48594 99200 48650 100000
rect 49422 99200 49478 100000
rect 50342 99200 50398 100000
rect 51262 99200 51318 100000
rect 52090 99200 52146 100000
rect 53010 99200 53066 100000
rect 53838 99200 53894 100000
rect 54758 99200 54814 100000
rect 55586 99200 55642 100000
rect 56506 99200 56562 100000
rect 57334 99200 57390 100000
rect 58254 99200 58310 100000
rect 59082 99200 59138 100000
rect 60002 99200 60058 100000
rect 60830 99200 60886 100000
rect 61750 99200 61806 100000
rect 62578 99200 62634 100000
rect 63498 99200 63554 100000
rect 64418 99200 64474 100000
rect 65246 99200 65302 100000
rect 66166 99200 66222 100000
rect 66994 99200 67050 100000
rect 67914 99200 67970 100000
rect 68742 99200 68798 100000
rect 69662 99200 69718 100000
rect 70490 99200 70546 100000
rect 71410 99200 71466 100000
rect 72238 99200 72294 100000
rect 73158 99200 73214 100000
rect 73986 99200 74042 100000
rect 74906 99200 74962 100000
rect 75826 99200 75882 100000
rect 76654 99200 76710 100000
rect 77574 99200 77630 100000
rect 78402 99200 78458 100000
rect 79322 99200 79378 100000
rect 80150 99200 80206 100000
rect 81070 99200 81126 100000
rect 81898 99200 81954 100000
rect 82818 99200 82874 100000
rect 83646 99200 83702 100000
rect 84566 99200 84622 100000
rect 85394 99200 85450 100000
rect 86314 99200 86370 100000
rect 87142 99200 87198 100000
rect 88062 99200 88118 100000
rect 88982 99200 89038 100000
rect 89810 99200 89866 100000
rect 90730 99200 90786 100000
rect 91558 99200 91614 100000
rect 92478 99200 92534 100000
rect 93306 99200 93362 100000
rect 94226 99200 94282 100000
rect 95054 99200 95110 100000
rect 95974 99200 96030 100000
rect 96802 99200 96858 100000
rect 97722 99200 97778 100000
rect 98550 99200 98606 100000
rect 99470 99200 99526 100000
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 662 0 718 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4526 0 4582 800
rect 4710 0 4766 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6366 0 6422 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17130 0 17186 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41602 0 41658 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43074 0 43130 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62946 0 63002 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64786 0 64842 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66626 0 66682 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70490 0 70546 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72882 0 72938 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74906 0 74962 800
rect 75090 0 75146 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78586 0 78642 800
rect 78770 0 78826 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82634 0 82690 800
rect 82818 0 82874 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86314 0 86370 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88706 0 88762 800
rect 88890 0 88946 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90546 0 90602 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92754 0 92810 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94410 0 94466 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96434 0 96490 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
<< obsm2 >>
rect 20 99144 330 99385
rect 498 99144 1158 99385
rect 1326 99144 2078 99385
rect 2246 99144 2906 99385
rect 3074 99144 3826 99385
rect 3994 99144 4654 99385
rect 4822 99144 5574 99385
rect 5742 99144 6402 99385
rect 6570 99144 7322 99385
rect 7490 99144 8150 99385
rect 8318 99144 9070 99385
rect 9238 99144 9898 99385
rect 10066 99144 10818 99385
rect 10986 99144 11646 99385
rect 11814 99144 12566 99385
rect 12734 99144 13486 99385
rect 13654 99144 14314 99385
rect 14482 99144 15234 99385
rect 15402 99144 16062 99385
rect 16230 99144 16982 99385
rect 17150 99144 17810 99385
rect 17978 99144 18730 99385
rect 18898 99144 19558 99385
rect 19726 99144 20478 99385
rect 20646 99144 21306 99385
rect 21474 99144 22226 99385
rect 22394 99144 23054 99385
rect 23222 99144 23974 99385
rect 24142 99144 24802 99385
rect 24970 99144 25722 99385
rect 25890 99144 26642 99385
rect 26810 99144 27470 99385
rect 27638 99144 28390 99385
rect 28558 99144 29218 99385
rect 29386 99144 30138 99385
rect 30306 99144 30966 99385
rect 31134 99144 31886 99385
rect 32054 99144 32714 99385
rect 32882 99144 33634 99385
rect 33802 99144 34462 99385
rect 34630 99144 35382 99385
rect 35550 99144 36210 99385
rect 36378 99144 37130 99385
rect 37298 99144 38050 99385
rect 38218 99144 38878 99385
rect 39046 99144 39798 99385
rect 39966 99144 40626 99385
rect 40794 99144 41546 99385
rect 41714 99144 42374 99385
rect 42542 99144 43294 99385
rect 43462 99144 44122 99385
rect 44290 99144 45042 99385
rect 45210 99144 45870 99385
rect 46038 99144 46790 99385
rect 46958 99144 47618 99385
rect 47786 99144 48538 99385
rect 48706 99144 49366 99385
rect 49534 99144 50286 99385
rect 50454 99144 51206 99385
rect 51374 99144 52034 99385
rect 52202 99144 52954 99385
rect 53122 99144 53782 99385
rect 53950 99144 54702 99385
rect 54870 99144 55530 99385
rect 55698 99144 56450 99385
rect 56618 99144 57278 99385
rect 57446 99144 58198 99385
rect 58366 99144 59026 99385
rect 59194 99144 59946 99385
rect 60114 99144 60774 99385
rect 60942 99144 61694 99385
rect 61862 99144 62522 99385
rect 62690 99144 63442 99385
rect 63610 99144 64362 99385
rect 64530 99144 65190 99385
rect 65358 99144 66110 99385
rect 66278 99144 66938 99385
rect 67106 99144 67858 99385
rect 68026 99144 68686 99385
rect 68854 99144 69606 99385
rect 69774 99144 70434 99385
rect 70602 99144 71354 99385
rect 71522 99144 72182 99385
rect 72350 99144 73102 99385
rect 73270 99144 73930 99385
rect 74098 99144 74850 99385
rect 75018 99144 75770 99385
rect 75938 99144 76598 99385
rect 76766 99144 77518 99385
rect 77686 99144 78346 99385
rect 78514 99144 79266 99385
rect 79434 99144 80094 99385
rect 80262 99144 81014 99385
rect 81182 99144 81842 99385
rect 82010 99144 82762 99385
rect 82930 99144 83590 99385
rect 83758 99144 84510 99385
rect 84678 99144 85338 99385
rect 85506 99144 86258 99385
rect 86426 99144 87086 99385
rect 87254 99144 88006 99385
rect 88174 99144 88926 99385
rect 89094 99144 89754 99385
rect 89922 99144 90674 99385
rect 90842 99144 91502 99385
rect 91670 99144 92422 99385
rect 92590 99144 93250 99385
rect 93418 99144 94170 99385
rect 94338 99144 94998 99385
rect 95166 99144 95918 99385
rect 96086 99144 96746 99385
rect 96914 99144 97666 99385
rect 97834 99144 98494 99385
rect 98662 99144 99414 99385
rect 99582 99144 99892 99385
rect 20 856 99892 99144
rect 20 575 54 856
rect 222 575 238 856
rect 406 575 422 856
rect 590 575 606 856
rect 774 575 790 856
rect 958 575 1066 856
rect 1234 575 1250 856
rect 1418 575 1434 856
rect 1602 575 1618 856
rect 1786 575 1802 856
rect 1970 575 2078 856
rect 2246 575 2262 856
rect 2430 575 2446 856
rect 2614 575 2630 856
rect 2798 575 2814 856
rect 2982 575 3090 856
rect 3258 575 3274 856
rect 3442 575 3458 856
rect 3626 575 3642 856
rect 3810 575 3826 856
rect 3994 575 4102 856
rect 4270 575 4286 856
rect 4454 575 4470 856
rect 4638 575 4654 856
rect 4822 575 4838 856
rect 5006 575 5114 856
rect 5282 575 5298 856
rect 5466 575 5482 856
rect 5650 575 5666 856
rect 5834 575 5850 856
rect 6018 575 6126 856
rect 6294 575 6310 856
rect 6478 575 6494 856
rect 6662 575 6678 856
rect 6846 575 6862 856
rect 7030 575 7138 856
rect 7306 575 7322 856
rect 7490 575 7506 856
rect 7674 575 7690 856
rect 7858 575 7874 856
rect 8042 575 8150 856
rect 8318 575 8334 856
rect 8502 575 8518 856
rect 8686 575 8702 856
rect 8870 575 8978 856
rect 9146 575 9162 856
rect 9330 575 9346 856
rect 9514 575 9530 856
rect 9698 575 9714 856
rect 9882 575 9990 856
rect 10158 575 10174 856
rect 10342 575 10358 856
rect 10526 575 10542 856
rect 10710 575 10726 856
rect 10894 575 11002 856
rect 11170 575 11186 856
rect 11354 575 11370 856
rect 11538 575 11554 856
rect 11722 575 11738 856
rect 11906 575 12014 856
rect 12182 575 12198 856
rect 12366 575 12382 856
rect 12550 575 12566 856
rect 12734 575 12750 856
rect 12918 575 13026 856
rect 13194 575 13210 856
rect 13378 575 13394 856
rect 13562 575 13578 856
rect 13746 575 13762 856
rect 13930 575 14038 856
rect 14206 575 14222 856
rect 14390 575 14406 856
rect 14574 575 14590 856
rect 14758 575 14774 856
rect 14942 575 15050 856
rect 15218 575 15234 856
rect 15402 575 15418 856
rect 15586 575 15602 856
rect 15770 575 15786 856
rect 15954 575 16062 856
rect 16230 575 16246 856
rect 16414 575 16430 856
rect 16598 575 16614 856
rect 16782 575 16890 856
rect 17058 575 17074 856
rect 17242 575 17258 856
rect 17426 575 17442 856
rect 17610 575 17626 856
rect 17794 575 17902 856
rect 18070 575 18086 856
rect 18254 575 18270 856
rect 18438 575 18454 856
rect 18622 575 18638 856
rect 18806 575 18914 856
rect 19082 575 19098 856
rect 19266 575 19282 856
rect 19450 575 19466 856
rect 19634 575 19650 856
rect 19818 575 19926 856
rect 20094 575 20110 856
rect 20278 575 20294 856
rect 20462 575 20478 856
rect 20646 575 20662 856
rect 20830 575 20938 856
rect 21106 575 21122 856
rect 21290 575 21306 856
rect 21474 575 21490 856
rect 21658 575 21674 856
rect 21842 575 21950 856
rect 22118 575 22134 856
rect 22302 575 22318 856
rect 22486 575 22502 856
rect 22670 575 22686 856
rect 22854 575 22962 856
rect 23130 575 23146 856
rect 23314 575 23330 856
rect 23498 575 23514 856
rect 23682 575 23698 856
rect 23866 575 23974 856
rect 24142 575 24158 856
rect 24326 575 24342 856
rect 24510 575 24526 856
rect 24694 575 24710 856
rect 24878 575 24986 856
rect 25154 575 25170 856
rect 25338 575 25354 856
rect 25522 575 25538 856
rect 25706 575 25814 856
rect 25982 575 25998 856
rect 26166 575 26182 856
rect 26350 575 26366 856
rect 26534 575 26550 856
rect 26718 575 26826 856
rect 26994 575 27010 856
rect 27178 575 27194 856
rect 27362 575 27378 856
rect 27546 575 27562 856
rect 27730 575 27838 856
rect 28006 575 28022 856
rect 28190 575 28206 856
rect 28374 575 28390 856
rect 28558 575 28574 856
rect 28742 575 28850 856
rect 29018 575 29034 856
rect 29202 575 29218 856
rect 29386 575 29402 856
rect 29570 575 29586 856
rect 29754 575 29862 856
rect 30030 575 30046 856
rect 30214 575 30230 856
rect 30398 575 30414 856
rect 30582 575 30598 856
rect 30766 575 30874 856
rect 31042 575 31058 856
rect 31226 575 31242 856
rect 31410 575 31426 856
rect 31594 575 31610 856
rect 31778 575 31886 856
rect 32054 575 32070 856
rect 32238 575 32254 856
rect 32422 575 32438 856
rect 32606 575 32622 856
rect 32790 575 32898 856
rect 33066 575 33082 856
rect 33250 575 33266 856
rect 33434 575 33450 856
rect 33618 575 33726 856
rect 33894 575 33910 856
rect 34078 575 34094 856
rect 34262 575 34278 856
rect 34446 575 34462 856
rect 34630 575 34738 856
rect 34906 575 34922 856
rect 35090 575 35106 856
rect 35274 575 35290 856
rect 35458 575 35474 856
rect 35642 575 35750 856
rect 35918 575 35934 856
rect 36102 575 36118 856
rect 36286 575 36302 856
rect 36470 575 36486 856
rect 36654 575 36762 856
rect 36930 575 36946 856
rect 37114 575 37130 856
rect 37298 575 37314 856
rect 37482 575 37498 856
rect 37666 575 37774 856
rect 37942 575 37958 856
rect 38126 575 38142 856
rect 38310 575 38326 856
rect 38494 575 38510 856
rect 38678 575 38786 856
rect 38954 575 38970 856
rect 39138 575 39154 856
rect 39322 575 39338 856
rect 39506 575 39522 856
rect 39690 575 39798 856
rect 39966 575 39982 856
rect 40150 575 40166 856
rect 40334 575 40350 856
rect 40518 575 40534 856
rect 40702 575 40810 856
rect 40978 575 40994 856
rect 41162 575 41178 856
rect 41346 575 41362 856
rect 41530 575 41546 856
rect 41714 575 41822 856
rect 41990 575 42006 856
rect 42174 575 42190 856
rect 42358 575 42374 856
rect 42542 575 42650 856
rect 42818 575 42834 856
rect 43002 575 43018 856
rect 43186 575 43202 856
rect 43370 575 43386 856
rect 43554 575 43662 856
rect 43830 575 43846 856
rect 44014 575 44030 856
rect 44198 575 44214 856
rect 44382 575 44398 856
rect 44566 575 44674 856
rect 44842 575 44858 856
rect 45026 575 45042 856
rect 45210 575 45226 856
rect 45394 575 45410 856
rect 45578 575 45686 856
rect 45854 575 45870 856
rect 46038 575 46054 856
rect 46222 575 46238 856
rect 46406 575 46422 856
rect 46590 575 46698 856
rect 46866 575 46882 856
rect 47050 575 47066 856
rect 47234 575 47250 856
rect 47418 575 47434 856
rect 47602 575 47710 856
rect 47878 575 47894 856
rect 48062 575 48078 856
rect 48246 575 48262 856
rect 48430 575 48446 856
rect 48614 575 48722 856
rect 48890 575 48906 856
rect 49074 575 49090 856
rect 49258 575 49274 856
rect 49442 575 49458 856
rect 49626 575 49734 856
rect 49902 575 49918 856
rect 50086 575 50102 856
rect 50270 575 50286 856
rect 50454 575 50562 856
rect 50730 575 50746 856
rect 50914 575 50930 856
rect 51098 575 51114 856
rect 51282 575 51298 856
rect 51466 575 51574 856
rect 51742 575 51758 856
rect 51926 575 51942 856
rect 52110 575 52126 856
rect 52294 575 52310 856
rect 52478 575 52586 856
rect 52754 575 52770 856
rect 52938 575 52954 856
rect 53122 575 53138 856
rect 53306 575 53322 856
rect 53490 575 53598 856
rect 53766 575 53782 856
rect 53950 575 53966 856
rect 54134 575 54150 856
rect 54318 575 54334 856
rect 54502 575 54610 856
rect 54778 575 54794 856
rect 54962 575 54978 856
rect 55146 575 55162 856
rect 55330 575 55346 856
rect 55514 575 55622 856
rect 55790 575 55806 856
rect 55974 575 55990 856
rect 56158 575 56174 856
rect 56342 575 56358 856
rect 56526 575 56634 856
rect 56802 575 56818 856
rect 56986 575 57002 856
rect 57170 575 57186 856
rect 57354 575 57370 856
rect 57538 575 57646 856
rect 57814 575 57830 856
rect 57998 575 58014 856
rect 58182 575 58198 856
rect 58366 575 58474 856
rect 58642 575 58658 856
rect 58826 575 58842 856
rect 59010 575 59026 856
rect 59194 575 59210 856
rect 59378 575 59486 856
rect 59654 575 59670 856
rect 59838 575 59854 856
rect 60022 575 60038 856
rect 60206 575 60222 856
rect 60390 575 60498 856
rect 60666 575 60682 856
rect 60850 575 60866 856
rect 61034 575 61050 856
rect 61218 575 61234 856
rect 61402 575 61510 856
rect 61678 575 61694 856
rect 61862 575 61878 856
rect 62046 575 62062 856
rect 62230 575 62246 856
rect 62414 575 62522 856
rect 62690 575 62706 856
rect 62874 575 62890 856
rect 63058 575 63074 856
rect 63242 575 63258 856
rect 63426 575 63534 856
rect 63702 575 63718 856
rect 63886 575 63902 856
rect 64070 575 64086 856
rect 64254 575 64270 856
rect 64438 575 64546 856
rect 64714 575 64730 856
rect 64898 575 64914 856
rect 65082 575 65098 856
rect 65266 575 65282 856
rect 65450 575 65558 856
rect 65726 575 65742 856
rect 65910 575 65926 856
rect 66094 575 66110 856
rect 66278 575 66294 856
rect 66462 575 66570 856
rect 66738 575 66754 856
rect 66922 575 66938 856
rect 67106 575 67122 856
rect 67290 575 67398 856
rect 67566 575 67582 856
rect 67750 575 67766 856
rect 67934 575 67950 856
rect 68118 575 68134 856
rect 68302 575 68410 856
rect 68578 575 68594 856
rect 68762 575 68778 856
rect 68946 575 68962 856
rect 69130 575 69146 856
rect 69314 575 69422 856
rect 69590 575 69606 856
rect 69774 575 69790 856
rect 69958 575 69974 856
rect 70142 575 70158 856
rect 70326 575 70434 856
rect 70602 575 70618 856
rect 70786 575 70802 856
rect 70970 575 70986 856
rect 71154 575 71170 856
rect 71338 575 71446 856
rect 71614 575 71630 856
rect 71798 575 71814 856
rect 71982 575 71998 856
rect 72166 575 72182 856
rect 72350 575 72458 856
rect 72626 575 72642 856
rect 72810 575 72826 856
rect 72994 575 73010 856
rect 73178 575 73194 856
rect 73362 575 73470 856
rect 73638 575 73654 856
rect 73822 575 73838 856
rect 74006 575 74022 856
rect 74190 575 74206 856
rect 74374 575 74482 856
rect 74650 575 74666 856
rect 74834 575 74850 856
rect 75018 575 75034 856
rect 75202 575 75310 856
rect 75478 575 75494 856
rect 75662 575 75678 856
rect 75846 575 75862 856
rect 76030 575 76046 856
rect 76214 575 76322 856
rect 76490 575 76506 856
rect 76674 575 76690 856
rect 76858 575 76874 856
rect 77042 575 77058 856
rect 77226 575 77334 856
rect 77502 575 77518 856
rect 77686 575 77702 856
rect 77870 575 77886 856
rect 78054 575 78070 856
rect 78238 575 78346 856
rect 78514 575 78530 856
rect 78698 575 78714 856
rect 78882 575 78898 856
rect 79066 575 79082 856
rect 79250 575 79358 856
rect 79526 575 79542 856
rect 79710 575 79726 856
rect 79894 575 79910 856
rect 80078 575 80094 856
rect 80262 575 80370 856
rect 80538 575 80554 856
rect 80722 575 80738 856
rect 80906 575 80922 856
rect 81090 575 81106 856
rect 81274 575 81382 856
rect 81550 575 81566 856
rect 81734 575 81750 856
rect 81918 575 81934 856
rect 82102 575 82118 856
rect 82286 575 82394 856
rect 82562 575 82578 856
rect 82746 575 82762 856
rect 82930 575 82946 856
rect 83114 575 83130 856
rect 83298 575 83406 856
rect 83574 575 83590 856
rect 83758 575 83774 856
rect 83942 575 83958 856
rect 84126 575 84234 856
rect 84402 575 84418 856
rect 84586 575 84602 856
rect 84770 575 84786 856
rect 84954 575 84970 856
rect 85138 575 85246 856
rect 85414 575 85430 856
rect 85598 575 85614 856
rect 85782 575 85798 856
rect 85966 575 85982 856
rect 86150 575 86258 856
rect 86426 575 86442 856
rect 86610 575 86626 856
rect 86794 575 86810 856
rect 86978 575 86994 856
rect 87162 575 87270 856
rect 87438 575 87454 856
rect 87622 575 87638 856
rect 87806 575 87822 856
rect 87990 575 88006 856
rect 88174 575 88282 856
rect 88450 575 88466 856
rect 88634 575 88650 856
rect 88818 575 88834 856
rect 89002 575 89018 856
rect 89186 575 89294 856
rect 89462 575 89478 856
rect 89646 575 89662 856
rect 89830 575 89846 856
rect 90014 575 90030 856
rect 90198 575 90306 856
rect 90474 575 90490 856
rect 90658 575 90674 856
rect 90842 575 90858 856
rect 91026 575 91042 856
rect 91210 575 91318 856
rect 91486 575 91502 856
rect 91670 575 91686 856
rect 91854 575 91870 856
rect 92038 575 92146 856
rect 92314 575 92330 856
rect 92498 575 92514 856
rect 92682 575 92698 856
rect 92866 575 92882 856
rect 93050 575 93158 856
rect 93326 575 93342 856
rect 93510 575 93526 856
rect 93694 575 93710 856
rect 93878 575 93894 856
rect 94062 575 94170 856
rect 94338 575 94354 856
rect 94522 575 94538 856
rect 94706 575 94722 856
rect 94890 575 94906 856
rect 95074 575 95182 856
rect 95350 575 95366 856
rect 95534 575 95550 856
rect 95718 575 95734 856
rect 95902 575 95918 856
rect 96086 575 96194 856
rect 96362 575 96378 856
rect 96546 575 96562 856
rect 96730 575 96746 856
rect 96914 575 96930 856
rect 97098 575 97206 856
rect 97374 575 97390 856
rect 97558 575 97574 856
rect 97742 575 97758 856
rect 97926 575 97942 856
rect 98110 575 98218 856
rect 98386 575 98402 856
rect 98570 575 98586 856
rect 98754 575 98770 856
rect 98938 575 98954 856
rect 99122 575 99230 856
rect 99398 575 99414 856
rect 99582 575 99598 856
rect 99766 575 99782 856
<< metal3 >>
rect 0 99288 800 99408
rect 0 98200 800 98320
rect 0 97112 800 97232
rect 0 96024 800 96144
rect 0 94936 800 95056
rect 0 93848 800 93968
rect 0 92760 800 92880
rect 0 91672 800 91792
rect 0 90584 800 90704
rect 0 89496 800 89616
rect 0 88408 800 88528
rect 0 87320 800 87440
rect 0 86232 800 86352
rect 0 85008 800 85128
rect 0 83920 800 84040
rect 0 82832 800 82952
rect 0 81744 800 81864
rect 0 80656 800 80776
rect 0 79568 800 79688
rect 0 78480 800 78600
rect 0 77392 800 77512
rect 0 76304 800 76424
rect 0 75216 800 75336
rect 0 74128 800 74248
rect 0 73040 800 73160
rect 0 71952 800 72072
rect 0 70728 800 70848
rect 0 69640 800 69760
rect 0 68552 800 68672
rect 0 67464 800 67584
rect 0 66376 800 66496
rect 0 65288 800 65408
rect 0 64200 800 64320
rect 0 63112 800 63232
rect 0 62024 800 62144
rect 0 60936 800 61056
rect 0 59848 800 59968
rect 0 58760 800 58880
rect 0 57672 800 57792
rect 0 56448 800 56568
rect 0 55360 800 55480
rect 0 54272 800 54392
rect 0 53184 800 53304
rect 0 52096 800 52216
rect 0 51008 800 51128
rect 0 49920 800 50040
rect 99200 49920 100000 50040
rect 0 48832 800 48952
rect 0 47744 800 47864
rect 0 46656 800 46776
rect 0 45568 800 45688
rect 0 44480 800 44600
rect 0 43392 800 43512
rect 0 42168 800 42288
rect 0 41080 800 41200
rect 0 39992 800 40112
rect 0 38904 800 39024
rect 0 37816 800 37936
rect 0 36728 800 36848
rect 0 35640 800 35760
rect 0 34552 800 34672
rect 0 33464 800 33584
rect 0 32376 800 32496
rect 0 31288 800 31408
rect 0 30200 800 30320
rect 0 29112 800 29232
rect 0 27888 800 28008
rect 0 26800 800 26920
rect 0 25712 800 25832
rect 0 24624 800 24744
rect 0 23536 800 23656
rect 0 22448 800 22568
rect 0 21360 800 21480
rect 0 20272 800 20392
rect 0 19184 800 19304
rect 0 18096 800 18216
rect 0 17008 800 17128
rect 0 15920 800 16040
rect 0 14832 800 14952
rect 0 13608 800 13728
rect 0 12520 800 12640
rect 0 11432 800 11552
rect 0 10344 800 10464
rect 0 9256 800 9376
rect 0 8168 800 8288
rect 0 7080 800 7200
rect 0 5992 800 6112
rect 0 4904 800 5024
rect 0 3816 800 3936
rect 0 2728 800 2848
rect 0 1640 800 1760
rect 0 552 800 672
<< obsm3 >>
rect 880 99208 99200 99381
rect 800 98400 99200 99208
rect 880 98120 99200 98400
rect 800 97312 99200 98120
rect 880 97032 99200 97312
rect 800 96224 99200 97032
rect 880 95944 99200 96224
rect 800 95136 99200 95944
rect 880 94856 99200 95136
rect 800 94048 99200 94856
rect 880 93768 99200 94048
rect 800 92960 99200 93768
rect 880 92680 99200 92960
rect 800 91872 99200 92680
rect 880 91592 99200 91872
rect 800 90784 99200 91592
rect 880 90504 99200 90784
rect 800 89696 99200 90504
rect 880 89416 99200 89696
rect 800 88608 99200 89416
rect 880 88328 99200 88608
rect 800 87520 99200 88328
rect 880 87240 99200 87520
rect 800 86432 99200 87240
rect 880 86152 99200 86432
rect 800 85208 99200 86152
rect 880 84928 99200 85208
rect 800 84120 99200 84928
rect 880 83840 99200 84120
rect 800 83032 99200 83840
rect 880 82752 99200 83032
rect 800 81944 99200 82752
rect 880 81664 99200 81944
rect 800 80856 99200 81664
rect 880 80576 99200 80856
rect 800 79768 99200 80576
rect 880 79488 99200 79768
rect 800 78680 99200 79488
rect 880 78400 99200 78680
rect 800 77592 99200 78400
rect 880 77312 99200 77592
rect 800 76504 99200 77312
rect 880 76224 99200 76504
rect 800 75416 99200 76224
rect 880 75136 99200 75416
rect 800 74328 99200 75136
rect 880 74048 99200 74328
rect 800 73240 99200 74048
rect 880 72960 99200 73240
rect 800 72152 99200 72960
rect 880 71872 99200 72152
rect 800 70928 99200 71872
rect 880 70648 99200 70928
rect 800 69840 99200 70648
rect 880 69560 99200 69840
rect 800 68752 99200 69560
rect 880 68472 99200 68752
rect 800 67664 99200 68472
rect 880 67384 99200 67664
rect 800 66576 99200 67384
rect 880 66296 99200 66576
rect 800 65488 99200 66296
rect 880 65208 99200 65488
rect 800 64400 99200 65208
rect 880 64120 99200 64400
rect 800 63312 99200 64120
rect 880 63032 99200 63312
rect 800 62224 99200 63032
rect 880 61944 99200 62224
rect 800 61136 99200 61944
rect 880 60856 99200 61136
rect 800 60048 99200 60856
rect 880 59768 99200 60048
rect 800 58960 99200 59768
rect 880 58680 99200 58960
rect 800 57872 99200 58680
rect 880 57592 99200 57872
rect 800 56648 99200 57592
rect 880 56368 99200 56648
rect 800 55560 99200 56368
rect 880 55280 99200 55560
rect 800 54472 99200 55280
rect 880 54192 99200 54472
rect 800 53384 99200 54192
rect 880 53104 99200 53384
rect 800 52296 99200 53104
rect 880 52016 99200 52296
rect 800 51208 99200 52016
rect 880 50928 99200 51208
rect 800 50120 99200 50928
rect 880 49840 99120 50120
rect 800 49032 99200 49840
rect 880 48752 99200 49032
rect 800 47944 99200 48752
rect 880 47664 99200 47944
rect 800 46856 99200 47664
rect 880 46576 99200 46856
rect 800 45768 99200 46576
rect 880 45488 99200 45768
rect 800 44680 99200 45488
rect 880 44400 99200 44680
rect 800 43592 99200 44400
rect 880 43312 99200 43592
rect 800 42368 99200 43312
rect 880 42088 99200 42368
rect 800 41280 99200 42088
rect 880 41000 99200 41280
rect 800 40192 99200 41000
rect 880 39912 99200 40192
rect 800 39104 99200 39912
rect 880 38824 99200 39104
rect 800 38016 99200 38824
rect 880 37736 99200 38016
rect 800 36928 99200 37736
rect 880 36648 99200 36928
rect 800 35840 99200 36648
rect 880 35560 99200 35840
rect 800 34752 99200 35560
rect 880 34472 99200 34752
rect 800 33664 99200 34472
rect 880 33384 99200 33664
rect 800 32576 99200 33384
rect 880 32296 99200 32576
rect 800 31488 99200 32296
rect 880 31208 99200 31488
rect 800 30400 99200 31208
rect 880 30120 99200 30400
rect 800 29312 99200 30120
rect 880 29032 99200 29312
rect 800 28088 99200 29032
rect 880 27808 99200 28088
rect 800 27000 99200 27808
rect 880 26720 99200 27000
rect 800 25912 99200 26720
rect 880 25632 99200 25912
rect 800 24824 99200 25632
rect 880 24544 99200 24824
rect 800 23736 99200 24544
rect 880 23456 99200 23736
rect 800 22648 99200 23456
rect 880 22368 99200 22648
rect 800 21560 99200 22368
rect 880 21280 99200 21560
rect 800 20472 99200 21280
rect 880 20192 99200 20472
rect 800 19384 99200 20192
rect 880 19104 99200 19384
rect 800 18296 99200 19104
rect 880 18016 99200 18296
rect 800 17208 99200 18016
rect 880 16928 99200 17208
rect 800 16120 99200 16928
rect 880 15840 99200 16120
rect 800 15032 99200 15840
rect 880 14752 99200 15032
rect 800 13808 99200 14752
rect 880 13528 99200 13808
rect 800 12720 99200 13528
rect 880 12440 99200 12720
rect 800 11632 99200 12440
rect 880 11352 99200 11632
rect 800 10544 99200 11352
rect 880 10264 99200 10544
rect 800 9456 99200 10264
rect 880 9176 99200 9456
rect 800 8368 99200 9176
rect 880 8088 99200 8368
rect 800 7280 99200 8088
rect 880 7000 99200 7280
rect 800 6192 99200 7000
rect 880 5912 99200 6192
rect 800 5104 99200 5912
rect 880 4824 99200 5104
rect 800 4016 99200 4824
rect 880 3736 99200 4016
rect 800 2928 99200 3736
rect 880 2648 99200 2928
rect 800 1840 99200 2648
rect 880 1560 99200 1840
rect 800 752 99200 1560
rect 880 579 99200 752
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 3187 2347 4128 84285
rect 4608 2347 19488 84285
rect 19968 2347 23861 84285
<< labels >>
rlabel metal2 s 386 99200 442 100000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 26698 99200 26754 100000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 29274 99200 29330 100000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 31942 99200 31998 100000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 34518 99200 34574 100000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 37186 99200 37242 100000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 39854 99200 39910 100000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 42430 99200 42486 100000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 45098 99200 45154 100000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47674 99200 47730 100000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 50342 99200 50398 100000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2962 99200 3018 100000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 53010 99200 53066 100000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 55586 99200 55642 100000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 58254 99200 58310 100000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 60830 99200 60886 100000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 63498 99200 63554 100000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 66166 99200 66222 100000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 68742 99200 68798 100000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 71410 99200 71466 100000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 73986 99200 74042 100000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 76654 99200 76710 100000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5630 99200 5686 100000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 79322 99200 79378 100000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 81898 99200 81954 100000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 84566 99200 84622 100000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 87142 99200 87198 100000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89810 99200 89866 100000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 92478 99200 92534 100000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 95054 99200 95110 100000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 97722 99200 97778 100000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8206 99200 8262 100000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10874 99200 10930 100000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13542 99200 13598 100000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16118 99200 16174 100000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18786 99200 18842 100000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 21362 99200 21418 100000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 24030 99200 24086 100000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 27526 99200 27582 100000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 30194 99200 30250 100000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32770 99200 32826 100000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 35438 99200 35494 100000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 38106 99200 38162 100000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 40682 99200 40738 100000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 43350 99200 43406 100000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 45926 99200 45982 100000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 48594 99200 48650 100000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 51262 99200 51318 100000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3882 99200 3938 100000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 53838 99200 53894 100000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 56506 99200 56562 100000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 59082 99200 59138 100000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 61750 99200 61806 100000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 64418 99200 64474 100000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66994 99200 67050 100000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 69662 99200 69718 100000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 72238 99200 72294 100000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 74906 99200 74962 100000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 77574 99200 77630 100000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6458 99200 6514 100000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 80150 99200 80206 100000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 82818 99200 82874 100000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 85394 99200 85450 100000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 88062 99200 88118 100000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 90730 99200 90786 100000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 93306 99200 93362 100000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 98550 99200 98606 100000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9126 99200 9182 100000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11702 99200 11758 100000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14370 99200 14426 100000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 17038 99200 17094 100000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19614 99200 19670 100000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 22282 99200 22338 100000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 24858 99200 24914 100000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2134 99200 2190 100000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 28446 99200 28502 100000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 31022 99200 31078 100000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 33690 99200 33746 100000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 36266 99200 36322 100000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 38934 99200 38990 100000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 41602 99200 41658 100000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 44178 99200 44234 100000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 46846 99200 46902 100000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 49422 99200 49478 100000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 52090 99200 52146 100000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 54758 99200 54814 100000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 57334 99200 57390 100000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 60002 99200 60058 100000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 62578 99200 62634 100000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 65246 99200 65302 100000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 67914 99200 67970 100000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 70490 99200 70546 100000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 73158 99200 73214 100000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 75826 99200 75882 100000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 78402 99200 78458 100000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7378 99200 7434 100000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 81070 99200 81126 100000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 83646 99200 83702 100000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 86314 99200 86370 100000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 88982 99200 89038 100000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 91558 99200 91614 100000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 94226 99200 94282 100000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 96802 99200 96858 100000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 99470 99200 99526 100000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9954 99200 10010 100000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12622 99200 12678 100000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15290 99200 15346 100000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 17866 99200 17922 100000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20534 99200 20590 100000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 23110 99200 23166 100000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 25778 99200 25834 100000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 ring0_clk
port 502 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 ring0_clkmux[0]
port 503 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 ring0_clkmux[1]
port 504 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 ring0_clkmux[2]
port 505 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 ring0_start
port 506 nsew signal output
rlabel metal3 s 0 552 800 672 6 ring0_trim_a[0]
port 507 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 ring0_trim_a[10]
port 508 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 ring0_trim_a[11]
port 509 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 ring0_trim_a[12]
port 510 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 ring0_trim_a[13]
port 511 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 ring0_trim_a[14]
port 512 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 ring0_trim_a[15]
port 513 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 ring0_trim_a[16]
port 514 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 ring0_trim_a[17]
port 515 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 ring0_trim_a[18]
port 516 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 ring0_trim_a[19]
port 517 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 ring0_trim_a[1]
port 518 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 ring0_trim_a[20]
port 519 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 ring0_trim_a[21]
port 520 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 ring0_trim_a[22]
port 521 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 ring0_trim_a[23]
port 522 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 ring0_trim_a[24]
port 523 nsew signal output
rlabel metal3 s 0 55360 800 55480 6 ring0_trim_a[25]
port 524 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 ring0_trim_a[26]
port 525 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 ring0_trim_a[27]
port 526 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 ring0_trim_a[2]
port 527 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 ring0_trim_a[3]
port 528 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 ring0_trim_a[4]
port 529 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 ring0_trim_a[5]
port 530 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 ring0_trim_a[6]
port 531 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 ring0_trim_a[7]
port 532 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 ring0_trim_a[8]
port 533 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 ring0_trim_a[9]
port 534 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 ring0_trim_b[0]
port 535 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 ring0_trim_b[10]
port 536 nsew signal output
rlabel metal3 s 0 71952 800 72072 6 ring0_trim_b[11]
port 537 nsew signal output
rlabel metal3 s 0 73040 800 73160 6 ring0_trim_b[12]
port 538 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 ring0_trim_b[13]
port 539 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 ring0_trim_b[14]
port 540 nsew signal output
rlabel metal3 s 0 76304 800 76424 6 ring0_trim_b[15]
port 541 nsew signal output
rlabel metal3 s 0 77392 800 77512 6 ring0_trim_b[16]
port 542 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 ring0_trim_b[17]
port 543 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 ring0_trim_b[18]
port 544 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 ring0_trim_b[19]
port 545 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 ring0_trim_b[1]
port 546 nsew signal output
rlabel metal3 s 0 81744 800 81864 6 ring0_trim_b[20]
port 547 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 ring0_trim_b[21]
port 548 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 ring0_trim_b[22]
port 549 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 ring0_trim_b[23]
port 550 nsew signal output
rlabel metal3 s 0 86232 800 86352 6 ring0_trim_b[24]
port 551 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 ring0_trim_b[25]
port 552 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 ring0_trim_b[26]
port 553 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 ring0_trim_b[27]
port 554 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 ring0_trim_b[2]
port 555 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 ring0_trim_b[3]
port 556 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 ring0_trim_b[4]
port 557 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 ring0_trim_b[5]
port 558 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 ring0_trim_b[6]
port 559 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 ring0_trim_b[7]
port 560 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 ring0_trim_b[8]
port 561 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 ring0_trim_b[9]
port 562 nsew signal output
rlabel metal3 s 99200 49920 100000 50040 6 ring1_clk
port 563 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 ring1_clkmux[0]
port 564 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 ring1_clkmux[1]
port 565 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 ring1_clkmux[2]
port 566 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 ring1_start
port 567 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 ring1_trim_a[0]
port 568 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 ring1_trim_a[10]
port 569 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 ring1_trim_a[11]
port 570 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 ring1_trim_a[12]
port 571 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 ring1_trim_a[13]
port 572 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 ring1_trim_a[14]
port 573 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 ring1_trim_a[15]
port 574 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 ring1_trim_a[16]
port 575 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 ring1_trim_a[17]
port 576 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 ring1_trim_a[18]
port 577 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 ring1_trim_a[19]
port 578 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 ring1_trim_a[1]
port 579 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 ring1_trim_a[20]
port 580 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 ring1_trim_a[21]
port 581 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 ring1_trim_a[22]
port 582 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 ring1_trim_a[23]
port 583 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 ring1_trim_a[24]
port 584 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 ring1_trim_a[25]
port 585 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 ring1_trim_a[2]
port 586 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 ring1_trim_a[3]
port 587 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 ring1_trim_a[4]
port 588 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 ring1_trim_a[5]
port 589 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 ring1_trim_a[6]
port 590 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 ring1_trim_a[7]
port 591 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 ring1_trim_a[8]
port 592 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 ring1_trim_a[9]
port 593 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 594 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 595 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 595 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 595 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 596 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 597 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 598 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[0]
port 599 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[10]
port 600 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[11]
port 601 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[12]
port 602 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[13]
port 603 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[14]
port 604 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[15]
port 605 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[16]
port 606 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[17]
port 607 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[18]
port 608 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[19]
port 609 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[1]
port 610 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[20]
port 611 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[21]
port 612 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[22]
port 613 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[23]
port 614 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[24]
port 615 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[25]
port 616 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[26]
port 617 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[27]
port 618 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[28]
port 619 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[29]
port 620 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[2]
port 621 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[30]
port 622 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[31]
port 623 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[3]
port 624 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[4]
port 625 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[5]
port 626 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[6]
port 627 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[7]
port 628 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[8]
port 629 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[9]
port 630 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_cyc_i
port 631 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[0]
port 632 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[10]
port 633 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[11]
port 634 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[12]
port 635 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[13]
port 636 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[14]
port 637 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[15]
port 638 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[16]
port 639 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[17]
port 640 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[18]
port 641 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[19]
port 642 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[1]
port 643 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[20]
port 644 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[21]
port 645 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[22]
port 646 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[23]
port 647 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[24]
port 648 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[25]
port 649 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[26]
port 650 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[27]
port 651 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[28]
port 652 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[29]
port 653 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[2]
port 654 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[30]
port 655 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[31]
port 656 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[3]
port 657 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[4]
port 658 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[5]
port 659 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[6]
port 660 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[7]
port 661 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[8]
port 662 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[9]
port 663 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_o[0]
port 664 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[10]
port 665 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[11]
port 666 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[12]
port 667 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[13]
port 668 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[14]
port 669 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[15]
port 670 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[16]
port 671 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[17]
port 672 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[18]
port 673 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[19]
port 674 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[1]
port 675 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[20]
port 676 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[21]
port 677 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[22]
port 678 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[23]
port 679 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[24]
port 680 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[25]
port 681 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[26]
port 682 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[27]
port 683 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[28]
port 684 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[29]
port 685 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_o[2]
port 686 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[30]
port 687 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[31]
port 688 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[3]
port 689 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[4]
port 690 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[5]
port 691 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_o[6]
port 692 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[7]
port 693 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[8]
port 694 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[9]
port 695 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_sel_i[0]
port 696 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[1]
port 697 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_sel_i[2]
port 698 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_sel_i[3]
port 699 nsew signal input
rlabel metal2 s 846 0 902 800 6 wbs_stb_i
port 700 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 701 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 100000 100000
string LEFview TRUE
string GDS_FILE /project/openlane/digitalcore_macro/runs/digitalcore_macro/results/magic/digitalcore_macro.gds
string GDS_END 9268786
string GDS_START 643032
<< end >>

